* SPICE NETLIST
***************************************

.SUBCKT nwell_contact
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT tri01 VDD GND
** N=8 EP=2 IP=2 FDC=6
M0 GND E 6 GND N L=4e-07 W=1e-06 AD=2.4e-12 AS=1.1e-12 $X=11500 $Y=31000 $D=1
M1 7 A GND GND N L=4e-07 W=2e-06 AD=1.2e-12 AS=2.4e-12 $X=20000 $Y=26000 $D=1
M2 Y E 7 GND N L=4e-07 W=2e-06 AD=2.2e-12 AS=1.2e-12 $X=25000 $Y=26000 $D=1
M3 VDD E 6 VDD P L=4e-07 W=1.8e-06 AD=4.32e-12 AS=1.58e-12 $X=11500 $Y=71000 $D=0
M4 8 A VDD VDD P L=4e-07 W=3.6e-06 AD=2.16e-12 AS=4.32e-12 $X=20000 $Y=71000 $D=0
M5 Y 6 8 VDD P L=4e-07 W=3.6e-06 AD=3.66e-12 AS=2.16e-12 $X=25000 $Y=71000 $D=0
.ENDS
***************************************
.SUBCKT nand02 GND
** N=6 EP=1 IP=2 FDC=4
M0 6 A1 GND GND N L=4e-07 W=2e-06 AD=1.2e-12 AS=2.2e-12 $X=11500 $Y=26000 $D=1
M1 Y A0 6 GND N L=4e-07 W=2e-06 AD=2.2e-12 AS=1.2e-12 $X=16500 $Y=26000 $D=1
M2 Y A1 VDD VDD P L=4e-07 W=2.4e-06 AD=2.88e-12 AS=2.44e-12 $X=11500 $Y=77000 $D=0
M3 VDD A0 Y VDD P L=4e-07 W=2.4e-06 AD=2.44e-12 AS=2.88e-12 $X=19500 $Y=77000 $D=0
.ENDS
***************************************
.SUBCKT oai22 GND VDD
** N=10 EP=2 IP=2 FDC=8
M0 Y A0 8 GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.2e-12 $X=11500 $Y=21000 $D=1
M1 8 A1 Y GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.4e-12 $X=19500 $Y=21000 $D=1
M2 GND B1 8 GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.4e-12 $X=27500 $Y=21000 $D=1
M3 8 B0 GND GND N L=4e-07 W=2e-06 AD=2.2e-12 AS=2.4e-12 $X=35500 $Y=21000 $D=1
M4 9 A0 VDD VDD P L=4e-07 W=4.8e-06 AD=2.88e-12 AS=4.88e-12 $X=15000 $Y=65000 $D=0
M5 Y A1 9 VDD P L=4e-07 W=4.8e-06 AD=5.76e-12 AS=2.88e-12 $X=20000 $Y=65000 $D=0
M6 10 B1 Y VDD P L=4e-07 W=4.8e-06 AD=2.88e-12 AS=5.76e-12 $X=28000 $Y=65000 $D=0
M7 VDD B0 10 VDD P L=4e-07 W=4.8e-06 AD=4.88e-12 AS=2.88e-12 $X=33000 $Y=65000 $D=0
.ENDS
***************************************
.SUBCKT inv02 GND VDD
** N=4 EP=2 IP=1 FDC=2
M0 Y A GND GND N L=4e-07 W=2e-06 AD=2.2e-12 AS=2.2e-12 $X=11500 $Y=26000 $D=1
M1 Y A VDD VDD P L=4e-07 W=3.6e-06 AD=3.66e-12 AS=3.66e-12 $X=11500 $Y=71000 $D=0
.ENDS
***************************************
.SUBCKT mux21_ni GND VDD
** N=12 EP=2 IP=0 FDC=12
M0 GND S0 7 GND N L=4e-07 W=1e-06 AD=2.4e-12 AS=1.1e-12 $X=11500 $Y=31000 $D=1
M1 9 S0 GND GND N L=4e-07 W=2e-06 AD=1.2e-12 AS=2.4e-12 $X=20000 $Y=26000 $D=1
M2 8 A1 9 GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=1.2e-12 $X=25000 $Y=26000 $D=1
M3 10 A0 8 GND N L=4e-07 W=2e-06 AD=1.2e-12 AS=2.4e-12 $X=33000 $Y=26000 $D=1
M4 GND 7 10 GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=1.2e-12 $X=38000 $Y=26000 $D=1
M5 Y 8 GND GND N L=4e-07 W=1e-06 AD=1.1e-12 AS=2.4e-12 $X=46500 $Y=31000 $D=1
M6 VDD S0 7 VDD P L=4e-07 W=1.8e-06 AD=4.32e-12 AS=1.58e-12 $X=11500 $Y=71000 $D=0
M7 11 S0 VDD VDD P L=4e-07 W=3.6e-06 AD=2.16e-12 AS=4.32e-12 $X=20000 $Y=71000 $D=0
M8 8 A0 11 VDD P L=4e-07 W=3.6e-06 AD=4.32e-12 AS=2.16e-12 $X=25000 $Y=71000 $D=0
M9 12 A1 8 VDD P L=4e-07 W=3.6e-06 AD=2.16e-12 AS=4.32e-12 $X=33000 $Y=71000 $D=0
M10 VDD 7 12 VDD P L=4e-07 W=3.6e-06 AD=4.32e-12 AS=2.16e-12 $X=38000 $Y=71000 $D=0
M11 Y 8 VDD VDD P L=4e-07 W=1.8e-06 AD=1.58e-12 AS=4.32e-12 $X=46500 $Y=71000 $D=0
.ENDS
***************************************
.SUBCKT mux21 GND VDD
** N=11 EP=2 IP=3 FDC=10
M0 8 7 Y GND N L=4e-07 W=2e-06 AD=1.2e-12 AS=2.2e-12 $X=11500 $Y=25000 $D=1
M1 GND A0 8 GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=1.2e-12 $X=16500 $Y=25000 $D=1
M2 9 A1 GND GND N L=4e-07 W=2e-06 AD=1.2e-12 AS=2.4e-12 $X=24500 $Y=25000 $D=1
M3 Y S0 9 GND N L=4e-07 W=2e-06 AD=2.2e-12 AS=1.2e-12 $X=29500 $Y=25000 $D=1
M4 GND S0 7 GND N L=4e-07 W=1e-06 AD=1.1e-12 AS=1.1e-12 $X=45500 $Y=30000 $D=1
M5 10 7 Y VDD P L=4e-07 W=3.6e-06 AD=2.16e-12 AS=3.66e-12 $X=13000 $Y=71000 $D=0
M6 VDD A1 10 VDD P L=4e-07 W=3.6e-06 AD=4.32e-12 AS=2.16e-12 $X=18000 $Y=71000 $D=0
M7 11 A0 VDD VDD P L=4e-07 W=3.6e-06 AD=2.16e-12 AS=4.32e-12 $X=26000 $Y=71000 $D=0
M8 Y S0 11 VDD P L=4e-07 W=3.6e-06 AD=3.66e-12 AS=2.16e-12 $X=31000 $Y=71000 $D=0
M9 VDD S0 7 VDD P L=4e-07 W=1.8e-06 AD=1.58e-12 AS=1.58e-12 $X=47000 $Y=71000 $D=0
.ENDS
***************************************
.SUBCKT dffr GND VDD
** N=23 EP=2 IP=9 FDC=34
M0 16 D GND GND N L=4e-07 W=3e-06 AD=1.8e-12 AS=3.3e-12 $X=11500 $Y=26000 $D=1
M1 8 12 16 GND N L=4e-07 W=3e-06 AD=3.5e-12 AS=1.8e-12 $X=16500 $Y=26000 $D=1
M2 17 11 8 GND N L=4e-07 W=1e-06 AD=6e-13 AS=3.5e-12 $X=25000 $Y=31000 $D=1
M3 GND 9 17 GND N L=4e-07 W=1e-06 AD=2.4e-12 AS=6e-13 $X=30000 $Y=31000 $D=1
M4 9 8 GND GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.4e-12 $X=38500 $Y=26000 $D=1
M5 GND R 9 GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.4e-12 $X=46500 $Y=26000 $D=1
M6 10 9 GND GND N L=4e-07 W=1e-06 AD=1.1e-12 AS=2.4e-12 $X=55000 $Y=31000 $D=1
M7 GND 12 11 GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.2e-12 $X=76000 $Y=31000 $D=1
M8 12 CLK GND GND N L=4e-07 W=2e-06 AD=2.2e-12 AS=2.4e-12 $X=84000 $Y=31000 $D=1
M9 18 10 GND GND N L=4e-07 W=3e-06 AD=1.8e-12 AS=3.3e-12 $X=100000 $Y=26000 $D=1
M10 13 11 18 GND N L=4e-07 W=3e-06 AD=3.5e-12 AS=1.8e-12 $X=105000 $Y=26000 $D=1
M11 14 12 13 GND N L=4e-07 W=1e-06 AD=1.1e-12 AS=3.5e-12 $X=113500 $Y=26000 $D=1
M12 14 R GND GND N L=4e-07 W=1e-06 AD=1.2e-12 AS=1.1e-12 $X=130500 $Y=26000 $D=1
M13 GND 15 14 GND N L=4e-07 W=1e-06 AD=1.2e-12 AS=1.2e-12 $X=138500 $Y=26000 $D=1
M14 15 13 GND GND N L=4e-07 W=1e-06 AD=1.1e-12 AS=1.2e-12 $X=146500 $Y=26000 $D=1
M15 GND 13 QB GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.2e-12 $X=162500 $Y=31000 $D=1
M16 Q QB GND GND N L=4e-07 W=2e-06 AD=2.2e-12 AS=2.4e-12 $X=170500 $Y=31000 $D=1
M17 19 11 VDD VDD P L=4e-07 W=5.4e-06 AD=3.24e-12 AS=5.74e-12 $X=11500 $Y=62000 $D=0
M18 8 D 19 VDD P L=4e-07 W=5.4e-06 AD=6.14e-12 AS=3.24e-12 $X=16500 $Y=62000 $D=0
M19 20 12 8 VDD P L=4e-07 W=1e-06 AD=6e-13 AS=6.14e-12 $X=25000 $Y=62000 $D=0
M20 VDD 9 20 VDD P L=4e-07 W=1e-06 AD=1.1e-12 AS=6e-13 $X=30000 $Y=62000 $D=0
M21 21 8 9 VDD P L=4e-07 W=2.4e-06 AD=1.44e-12 AS=2.44e-12 $X=46000 $Y=62000 $D=0
M22 VDD R 21 VDD P L=4e-07 W=2.4e-06 AD=3e-12 AS=1.44e-12 $X=51000 $Y=62000 $D=0
M23 10 9 VDD VDD P L=4e-07 W=1.8e-06 AD=1.58e-12 AS=3e-12 $X=59500 $Y=62000 $D=0
M24 VDD 12 11 VDD P L=4e-07 W=3.6e-06 AD=4.32e-12 AS=3.66e-12 $X=76000 $Y=62000 $D=0
M25 12 CLK VDD VDD P L=4e-07 W=3.6e-06 AD=3.66e-12 AS=4.32e-12 $X=84000 $Y=62000 $D=0
M26 22 10 VDD VDD P L=4e-07 W=5.4e-06 AD=3.24e-12 AS=5.74e-12 $X=100000 $Y=53000 $D=0
M27 13 12 22 VDD P L=4e-07 W=5.4e-06 AD=6.14e-12 AS=3.24e-12 $X=105000 $Y=53000 $D=0
M28 14 11 13 VDD P L=4e-07 W=1e-06 AD=1.2e-12 AS=6.14e-12 $X=113500 $Y=68000 $D=0
M29 23 R 14 VDD P L=4e-07 W=1e-06 AD=6e-13 AS=1.2e-12 $X=121500 $Y=68000 $D=0
M30 VDD 15 23 VDD P L=4e-07 W=1e-06 AD=1.2e-12 AS=6e-13 $X=126500 $Y=68000 $D=0
M31 15 13 VDD VDD P L=4e-07 W=1e-06 AD=1.1e-12 AS=1.2e-12 $X=134500 $Y=68000 $D=0
M32 VDD 13 QB VDD P L=4e-07 W=3.6e-06 AD=4.32e-12 AS=3.66e-12 $X=162500 $Y=62000 $D=0
M33 Q QB VDD VDD P L=4e-07 W=3.6e-06 AD=3.66e-12 AS=4.32e-12 $X=170500 $Y=62000 $D=0
.ENDS
***************************************
.SUBCKT inv01 GND VDD
** N=4 EP=2 IP=1 FDC=2
M0 Y A GND GND N L=4e-07 W=1e-06 AD=1.1e-12 AS=1.1e-12 $X=11500 $Y=26000 $D=1
M1 Y A VDD VDD P L=4e-07 W=1.8e-06 AD=1.58e-12 AS=1.58e-12 $X=11500 $Y=80000 $D=0
.ENDS
***************************************
.SUBCKT buf02 GND VDD
** N=5 EP=2 IP=1 FDC=4
M0 GND 5 Y GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.2e-12 $X=11500 $Y=26000 $D=1
M1 5 A GND GND N L=4e-07 W=1e-06 AD=1.1e-12 AS=2.4e-12 $X=20000 $Y=31000 $D=1
M2 VDD 5 Y VDD P L=4e-07 W=3.6e-06 AD=4.32e-12 AS=3.66e-12 $X=11500 $Y=71000 $D=0
M3 5 A VDD VDD P L=4e-07 W=1.8e-06 AD=1.58e-12 AS=4.32e-12 $X=20000 $Y=71000 $D=0
.ENDS
***************************************
.SUBCKT aoi22 VDD GND
** N=10 EP=2 IP=2 FDC=8
M0 9 B1 GND GND N L=4e-07 W=2e-06 AD=1.2e-12 AS=2.2e-12 $X=14500 $Y=26000 $D=1
M1 Y B0 9 GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=1.2e-12 $X=19500 $Y=26000 $D=1
M2 10 A0 Y GND N L=4e-07 W=2e-06 AD=1.2e-12 AS=2.4e-12 $X=27500 $Y=26000 $D=1
M3 GND A1 10 GND N L=4e-07 W=2e-06 AD=2.2e-12 AS=1.2e-12 $X=32500 $Y=26000 $D=1
M4 Y B1 8 VDD P L=4e-07 W=2.6e-06 AD=3.12e-12 AS=2.56e-12 $X=11500 $Y=76000 $D=0
M5 8 B0 Y VDD P L=4e-07 W=2.6e-06 AD=3.12e-12 AS=3.12e-12 $X=19500 $Y=76000 $D=0
M6 VDD A0 8 VDD P L=4e-07 W=2.6e-06 AD=3.12e-12 AS=3.12e-12 $X=27500 $Y=76000 $D=0
M7 8 A1 VDD VDD P L=4e-07 W=2.6e-06 AD=2.56e-12 AS=3.12e-12 $X=35500 $Y=76000 $D=0
.ENDS
***************************************
.SUBCKT ICV_1 1 2
** N=2 EP=2 IP=4 FDC=46
X0 1 2 mux21_ni $T=-60000 0 0 0 $X=-60000 $Y=0
X1 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_2 1 2
** N=2 EP=2 IP=4 FDC=68
X0 1 2 dffr $T=-184000 0 0 0 $X=-184000 $Y=0
X1 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_3 1
** N=2 EP=1 IP=4 FDC=40
X0 2 1 tri01 $T=184000 0 0 0 $X=184000 $Y=0
X1 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_4 1 2
** N=2 EP=2 IP=4 FDC=68
X0 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
X1 1 2 dffr $T=184000 0 0 0 $X=184000 $Y=0
.ENDS
***************************************
.SUBCKT nand04 GND VDD
** N=10 EP=2 IP=2 FDC=8
M0 8 A0 Y GND N L=4e-07 W=4e-06 AD=2.4e-12 AS=4.4e-12 $X=11500 $Y=28000 $D=1
M1 9 A1 8 GND N L=4e-07 W=4e-06 AD=2.4e-12 AS=2.4e-12 $X=16500 $Y=28000 $D=1
M2 10 A2 9 GND N L=4e-07 W=4e-06 AD=2.4e-12 AS=2.4e-12 $X=21500 $Y=28000 $D=1
M3 GND A3 10 GND N L=4e-07 W=4e-06 AD=4.4e-12 AS=2.4e-12 $X=26500 $Y=28000 $D=1
M4 Y A0 VDD VDD P L=4e-07 W=4e-06 AD=4.8e-12 AS=4.4e-12 $X=11500 $Y=79500 $D=0
M5 VDD A1 Y VDD P L=4e-07 W=4e-06 AD=4.8e-12 AS=4.8e-12 $X=19500 $Y=79500 $D=0
M6 Y A2 VDD VDD P L=4e-07 W=4e-06 AD=4.8e-12 AS=4.8e-12 $X=27500 $Y=79500 $D=0
M7 VDD A3 Y VDD P L=4e-07 W=4e-06 AD=4.4e-12 AS=4.8e-12 $X=35500 $Y=79500 $D=0
.ENDS
***************************************
.SUBCKT oai221 GND
** N=12 EP=1 IP=3 FDC=10
M0 8 C0 GND GND N L=4e-07 W=3e-06 AD=3.3e-12 AS=3.3e-12 $X=11500 $Y=25000 $D=1
M1 Y A0 10 GND N L=4e-07 W=3e-06 AD=3.6e-12 AS=3.3e-12 $X=28000 $Y=25000 $D=1
M2 10 A1 Y GND N L=4e-07 W=3e-06 AD=3.6e-12 AS=3.6e-12 $X=36000 $Y=25000 $D=1
M3 8 B1 10 GND N L=4e-07 W=3e-06 AD=3.6e-12 AS=3.6e-12 $X=44000 $Y=25000 $D=1
M4 10 B0 8 GND N L=4e-07 W=3e-06 AD=3.3e-12 AS=3.6e-12 $X=52000 $Y=25000 $D=1
M5 VDD C0 Y VDD P L=4e-07 W=3e-06 AD=7.2e-12 AS=3.3e-12 $X=19500 $Y=74000 $D=0
M6 11 A0 VDD VDD P L=4e-07 W=6e-06 AD=3.6e-12 AS=7.2e-12 $X=28000 $Y=74000 $D=0
M7 Y A1 11 VDD P L=4e-07 W=6e-06 AD=7.2e-12 AS=3.6e-12 $X=33000 $Y=74000 $D=0
M8 12 B1 Y VDD P L=4e-07 W=6e-06 AD=3.6e-12 AS=7.2e-12 $X=41000 $Y=74000 $D=0
M9 VDD B0 12 VDD P L=4e-07 W=6e-06 AD=6.6e-12 AS=3.6e-12 $X=46000 $Y=74000 $D=0
.ENDS
***************************************
.SUBCKT ICV_5 1
** N=2 EP=1 IP=4 FDC=46
X0 1 2 mux21_ni $T=0 0 1 180 $X=-60000 $Y=0
X1 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_6 1 2
** N=2 EP=2 IP=4 FDC=46
X0 1 2 mux21_ni $T=184000 0 0 0 $X=184000 $Y=0
X1 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_7 1 2
** N=2 EP=2 IP=4 FDC=68
X0 1 2 dffr $T=0 0 1 180 $X=-184000 $Y=0
X1 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_8 1
** N=2 EP=1 IP=4 FDC=38
X0 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
X1 1 2 buf02 $T=217500 0 1 180 $X=184000 $Y=0
.ENDS
***************************************
.SUBCKT ICV_9 1 2
** N=2 EP=2 IP=4 FDC=42
X0 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
X1 2 1 aoi22 $T=184000 0 0 0 $X=184000 $Y=0
.ENDS
***************************************
.SUBCKT dff GND VDD
** N=20 EP=2 IP=5 FDC=28
M0 13 9 7 GND N L=4e-07 W=3e-06 AD=1.8e-12 AS=3.3e-12 $X=11500 $Y=26000 $D=1
M1 GND D 13 GND N L=4e-07 W=3e-06 AD=3.3e-12 AS=1.8e-12 $X=16500 $Y=26000 $D=1
M2 14 10 7 GND N L=4e-07 W=1e-06 AD=6e-13 AS=1.1e-12 $X=32500 $Y=36000 $D=1
M3 GND 8 14 GND N L=4e-07 W=1e-06 AD=1.2e-12 AS=6e-13 $X=37500 $Y=36000 $D=1
M4 8 7 GND GND N L=4e-07 W=1e-06 AD=1.1e-12 AS=1.2e-12 $X=45500 $Y=36000 $D=1
M5 GND CLK 9 GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.2e-12 $X=61500 $Y=28500 $D=1
M6 10 9 GND GND N L=4e-07 W=2e-06 AD=2.2e-12 AS=2.4e-12 $X=69500 $Y=28500 $D=1
M7 GND 12 11 GND N L=4e-07 W=1e-06 AD=1.2e-12 AS=1.1e-12 $X=85500 $Y=37500 $D=1
M8 15 11 GND GND N L=4e-07 W=1e-06 AD=6e-13 AS=1.2e-12 $X=93500 $Y=37500 $D=1
M9 12 9 15 GND N L=4e-07 W=1e-06 AD=1.1e-12 AS=6e-13 $X=98500 $Y=37500 $D=1
M10 16 7 GND GND N L=4e-07 W=3e-06 AD=1.8e-12 AS=3.3e-12 $X=115500 $Y=27500 $D=1
M11 12 10 16 GND N L=4e-07 W=3e-06 AD=3.3e-12 AS=1.8e-12 $X=120500 $Y=27500 $D=1
M12 GND 12 QB GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.2e-12 $X=136500 $Y=32500 $D=1
M13 Q QB GND GND N L=4e-07 W=2e-06 AD=2.2e-12 AS=2.4e-12 $X=144500 $Y=32500 $D=1
M14 17 D VDD VDD P L=4e-07 W=5.4e-06 AD=3.24e-12 AS=5.74e-12 $X=11500 $Y=62000 $D=0
M15 7 10 17 VDD P L=4e-07 W=5.4e-06 AD=6.14e-12 AS=3.24e-12 $X=16500 $Y=62000 $D=0
M16 18 9 7 VDD P L=4e-07 W=1e-06 AD=3.1e-12 AS=6.14e-12 $X=25000 $Y=84000 $D=0
M17 VDD 8 18 VDD P L=4e-07 W=1e-06 AD=1.2e-12 AS=3.1e-12 $X=32000 $Y=66500 $D=0
M18 8 7 VDD VDD P L=4e-07 W=1e-06 AD=1.1e-12 AS=1.2e-12 $X=40000 $Y=66500 $D=0
M19 VDD CLK 9 VDD P L=4e-07 W=3.6e-06 AD=4.32e-12 AS=3.66e-12 $X=61500 $Y=71000 $D=0
M20 10 9 VDD VDD P L=4e-07 W=3.6e-06 AD=3.66e-12 AS=4.32e-12 $X=69500 $Y=71000 $D=0
M21 VDD 12 11 VDD P L=4e-07 W=1e-06 AD=1.2e-12 AS=1.1e-12 $X=85500 $Y=84000 $D=0
M22 19 11 VDD VDD P L=4e-07 W=1e-06 AD=6e-13 AS=1.2e-12 $X=93500 $Y=84000 $D=0
M23 12 10 19 VDD P L=4e-07 W=1e-06 AD=6.14e-12 AS=6e-13 $X=98500 $Y=84000 $D=0
M24 20 9 12 VDD P L=4e-07 W=5.4e-06 AD=3.24e-12 AS=6.14e-12 $X=107000 $Y=62000 $D=0
M25 VDD 7 20 VDD P L=4e-07 W=5.4e-06 AD=5.74e-12 AS=3.24e-12 $X=112000 $Y=62000 $D=0
M26 VDD 12 QB VDD P L=4e-07 W=3.6e-06 AD=4.32e-12 AS=3.66e-12 $X=136500 $Y=71000 $D=0
M27 Q QB VDD VDD P L=4e-07 W=3.6e-06 AD=3.66e-12 AS=4.32e-12 $X=144500 $Y=71000 $D=0
.ENDS
***************************************
.SUBCKT ICV_10 1
** N=2 EP=1 IP=4 FDC=42
X0 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
X1 1 2 nand04 $T=184000 0 0 0 $X=184000 $Y=0
.ENDS
***************************************
.SUBCKT and03 GND VDD
** N=9 EP=2 IP=2 FDC=8
M0 8 A0 7 GND N L=4e-07 W=3e-06 AD=1.8e-12 AS=3.3e-12 $X=15500 $Y=18500 $D=1
M1 9 A1 8 GND N L=4e-07 W=3e-06 AD=1.8e-12 AS=1.8e-12 $X=20500 $Y=18500 $D=1
M2 GND A2 9 GND N L=4e-07 W=3e-06 AD=3.5e-12 AS=1.8e-12 $X=25500 $Y=18500 $D=1
M3 Y 7 GND GND N L=4e-07 W=1e-06 AD=1.1e-12 AS=3.5e-12 $X=34000 $Y=18500 $D=1
M4 VDD 7 Y VDD P L=4e-07 W=1.8e-06 AD=3.66e-12 AS=1.58e-12 $X=11500 $Y=86000 $D=0
M5 7 A0 VDD VDD P L=4e-07 W=3e-06 AD=3.6e-12 AS=3.66e-12 $X=20000 $Y=86000 $D=0
M6 VDD A1 7 VDD P L=4e-07 W=3e-06 AD=3.6e-12 AS=3.6e-12 $X=28000 $Y=86000 $D=0
M7 7 A2 VDD VDD P L=4e-07 W=3e-06 AD=3.3e-12 AS=3.6e-12 $X=36000 $Y=86000 $D=0
.ENDS
***************************************
.SUBCKT ICV_11 1 2
** N=2 EP=2 IP=4 FDC=80
X0 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
X1 1 2 ICV_1 $T=368000 0 1 180 $X=184000 $Y=0
.ENDS
***************************************
.SUBCKT ICV_12 1
** N=2 EP=1 IP=4 FDC=38
X0 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
X1 1 2 buf02 $T=184000 0 0 0 $X=184000 $Y=0
.ENDS
***************************************
.SUBCKT ICV_13 1 2
** N=2 EP=2 IP=4 FDC=36
X0 1 2 inv02 $T=184000 0 0 0 $X=184000 $Y=0
X1 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_14 1
** N=2 EP=1 IP=4 FDC=42
X0 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
X1 2 1 aoi22 $T=0 0 1 180 $X=-49000 $Y=0
.ENDS
***************************************
.SUBCKT ICV_15 1
** N=2 EP=1 IP=4 FDC=80
X0 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
X1 1 2 ICV_1 $T=-184000 0 0 0 $X=-244000 $Y=0
.ENDS
***************************************
.SUBCKT ICV_16 1 2
** N=2 EP=2 IP=4 FDC=42
X0 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
X1 2 1 aoi22 $T=233000 0 1 180 $X=184000 $Y=0
.ENDS
***************************************
.SUBCKT ICV_17 1 2
** N=2 EP=2 IP=4 FDC=68
X0 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
X1 1 2 dffr $T=368000 0 1 180 $X=184000 $Y=0
.ENDS
***************************************
.SUBCKT xnor2 GND VDD
** N=9 EP=2 IP=3 FDC=10
M0 7 6 GND GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.2e-12 $X=11500 $Y=26000 $D=1
M1 Y A0 7 GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.4e-12 $X=19500 $Y=26000 $D=1
M2 7 A1 Y GND N L=4e-07 W=2e-06 AD=2.2e-12 AS=2.4e-12 $X=27500 $Y=26000 $D=1
M3 8 A1 GND GND N L=4e-07 W=2e-06 AD=1.2e-12 AS=2.2e-12 $X=44500 $Y=26000 $D=1
M4 6 A0 8 GND N L=4e-07 W=2e-06 AD=2.2e-12 AS=1.2e-12 $X=49500 $Y=26000 $D=1
M5 VDD 6 Y VDD P L=4e-07 W=2.6e-06 AD=3.12e-12 AS=2.56e-12 $X=11500 $Y=76000 $D=0
M6 6 A0 VDD VDD P L=4e-07 W=2.6e-06 AD=3.12e-12 AS=3.12e-12 $X=19500 $Y=76000 $D=0
M7 VDD A1 6 VDD P L=4e-07 W=2.6e-06 AD=2.56e-12 AS=3.12e-12 $X=27500 $Y=76000 $D=0
M8 9 A1 Y VDD P L=4e-07 W=5.2e-06 AD=3.12e-12 AS=5.62e-12 $X=44500 $Y=63000 $D=0
M9 VDD A0 9 VDD P L=4e-07 W=5.2e-06 AD=5.62e-12 AS=3.12e-12 $X=49500 $Y=63000 $D=0
.ENDS
***************************************
.SUBCKT ICV_18 1 2
** N=3 EP=2 IP=4 FDC=22
X0 1 3 mux21_ni $T=64000 0 0 0 $X=64000 $Y=0
X1 1 2 xnor2 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT xor2 GND
** N=10 EP=1 IP=3 FDC=12
M0 9 A0 5 GND N L=4e-07 W=2e-06 AD=1.2e-12 AS=2.2e-12 $X=11500 $Y=26000 $D=1
M1 GND A1 9 GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=1.2e-12 $X=16500 $Y=26000 $D=1
M2 6 5 GND GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.4e-12 $X=24500 $Y=26000 $D=1
M3 8 A0 6 GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.4e-12 $X=32500 $Y=26000 $D=1
M4 6 A1 8 GND N L=4e-07 W=2e-06 AD=2.2e-12 AS=2.4e-12 $X=40500 $Y=26000 $D=1
M5 Y 8 GND GND N L=4e-07 W=1e-06 AD=1.1e-12 AS=1.1e-12 $X=56500 $Y=31000 $D=1
M6 5 A0 VDD VDD P L=4e-07 W=2.6e-06 AD=6.12e-12 AS=2.56e-12 $X=14500 $Y=63000 $D=0
M7 VDD A1 5 VDD P L=4e-07 W=2.6e-06 AD=6.14e-12 AS=6.12e-12 $X=23500 $Y=76000 $D=0
M8 10 A0 VDD VDD P L=4e-07 W=5.2e-06 AD=3.12e-12 AS=6.14e-12 $X=32000 $Y=63000 $D=0
M9 8 A1 10 VDD P L=4e-07 W=5.2e-06 AD=6.14e-12 AS=3.12e-12 $X=37000 $Y=63000 $D=0
M10 VDD 5 8 VDD P L=4e-07 W=2.6e-06 AD=3.22e-12 AS=6.14e-12 $X=45500 $Y=63000 $D=0
M11 Y 8 VDD VDD P L=4e-07 W=1.8e-06 AD=1.58e-12 AS=3.22e-12 $X=54000 $Y=63000 $D=0
.ENDS
***************************************
.SUBCKT ICV_19 1 2
** N=2 EP=2 IP=4 FDC=46
X0 1 2 mux21_ni $T=244000 0 1 180 $X=184000 $Y=0
X1 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_20 1
** N=3 EP=1 IP=4 FDC=20
X0 1 2 xnor2 $T=0 0 0 0 $X=0 $Y=0
X1 1 3 xnor2 $T=64000 0 0 0 $X=64000 $Y=0
.ENDS
***************************************
.SUBCKT ICV_21 1
** N=2 EP=1 IP=4 FDC=36
X0 1 2 inv02 $T=-25000 0 0 0 $X=-25000 $Y=0
X1 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_22 1
** N=3 EP=1 IP=4 FDC=18
X0 1 2 oai22 $T=-50000 0 0 0 $X=-50000 $Y=0
X1 1 3 xnor2 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_23 1 2
** N=2 EP=2 IP=4 FDC=42
X0 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
X1 1 2 and03 $T=184000 0 0 0 $X=184000 $Y=0
.ENDS
***************************************
.SUBCKT ICV_24 1
** N=2 EP=1 IP=4 FDC=80
X0 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
X1 1 2 ICV_6 $T=184000 0 0 0 $X=184000 $Y=0
.ENDS
***************************************
.SUBCKT ICV_25 1
** N=3 EP=1 IP=4 FDC=18
X0 2 1 aoi22 $T=113000 0 1 180 $X=64000 $Y=0
X1 1 3 xnor2 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT oai32 GND
** N=12 EP=1 IP=3 FDC=10
M0 9 A0 Y GND N L=4e-07 W=3e-06 AD=3.6e-12 AS=3.3e-12 $X=11500 $Y=18500 $D=1
M1 Y A1 9 GND N L=4e-07 W=3e-06 AD=3.6e-12 AS=3.6e-12 $X=19500 $Y=18500 $D=1
M2 9 A2 Y GND N L=4e-07 W=3e-06 AD=3.6e-12 AS=3.6e-12 $X=27500 $Y=18500 $D=1
M3 GND B1 9 GND N L=4e-07 W=3e-06 AD=3.6e-12 AS=3.6e-12 $X=35500 $Y=18500 $D=1
M4 9 B0 GND GND N L=4e-07 W=3e-06 AD=3.3e-12 AS=3.6e-12 $X=43500 $Y=18500 $D=1
M5 10 A0 VDD VDD P L=4e-07 W=7.2e-06 AD=4.32e-12 AS=7.82e-12 $X=16000 $Y=68000 $D=0
M6 11 A1 10 VDD P L=4e-07 W=7.2e-06 AD=4.32e-12 AS=4.32e-12 $X=21000 $Y=68000 $D=0
M7 Y A2 11 VDD P L=4e-07 W=7.2e-06 AD=8.88e-12 AS=4.32e-12 $X=26000 $Y=68000 $D=0
M8 12 B1 Y VDD P L=4e-07 W=4.8e-06 AD=2.88e-12 AS=8.88e-12 $X=34500 $Y=68000 $D=0
M9 VDD B0 12 VDD P L=4e-07 W=4.8e-06 AD=4.88e-12 AS=2.88e-12 $X=39500 $Y=68000 $D=0
.ENDS
***************************************
.SUBCKT or04 GND
** N=11 EP=1 IP=3 FDC=10
M0 GND 8 Y GND N L=4e-07 W=1e-06 AD=1.1e-12 AS=1.1e-12 $X=11500 $Y=26000 $D=1
M1 GND A0 8 GND N L=4e-07 W=1e-06 AD=1.2e-12 AS=1.1e-12 $X=27500 $Y=26000 $D=1
M2 8 A1 GND GND N L=4e-07 W=1e-06 AD=1.2e-12 AS=1.2e-12 $X=35500 $Y=26000 $D=1
M3 GND A2 8 GND N L=4e-07 W=1e-06 AD=1.2e-12 AS=1.2e-12 $X=43500 $Y=26000 $D=1
M4 8 A3 GND GND N L=4e-07 W=1e-06 AD=1.1e-12 AS=1.2e-12 $X=51500 $Y=26000 $D=1
M5 VDD 8 Y VDD P L=4e-07 W=1.8e-06 AD=4.32e-12 AS=1.58e-12 $X=23500 $Y=71000 $D=0
M6 9 A0 VDD VDD P L=4e-07 W=3.6e-06 AD=2.16e-12 AS=4.32e-12 $X=32000 $Y=71000 $D=0
M7 10 A1 9 VDD P L=4e-07 W=3.6e-06 AD=2.16e-12 AS=2.16e-12 $X=37000 $Y=71000 $D=0
M8 11 A2 10 VDD P L=4e-07 W=3.6e-06 AD=2.16e-12 AS=2.16e-12 $X=42000 $Y=71000 $D=0
M9 8 A3 11 VDD P L=4e-07 W=3.6e-06 AD=3.66e-12 AS=2.16e-12 $X=47000 $Y=71000 $D=0
.ENDS
***************************************
.SUBCKT and02 GND VDD
** N=7 EP=2 IP=2 FDC=6
M0 7 A0 6 GND N L=4e-07 W=2e-06 AD=1.2e-12 AS=2.2e-12 $X=14500 $Y=26000 $D=1
M1 GND A1 7 GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=1.2e-12 $X=19500 $Y=26000 $D=1
M2 Y 6 GND GND N L=4e-07 W=1e-06 AD=1.1e-12 AS=2.4e-12 $X=28000 $Y=31000 $D=1
M3 6 A0 VDD VDD P L=4e-07 W=2.4e-06 AD=2.88e-12 AS=2.44e-12 $X=11500 $Y=77000 $D=0
M4 VDD A1 6 VDD P L=4e-07 W=2.4e-06 AD=3e-12 AS=2.88e-12 $X=19500 $Y=77000 $D=0
M5 Y 6 VDD VDD P L=4e-07 W=1.8e-06 AD=1.58e-12 AS=3e-12 $X=28000 $Y=77000 $D=0
.ENDS
***************************************
.SUBCKT ICV_26 1
** N=2 EP=1 IP=4 FDC=36
X0 1 2 inv02 $T=209000 0 1 180 $X=184000 $Y=0
X1 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT nor02_2x GND
** N=6 EP=1 IP=0 FDC=4
M0 Y A0 GND GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.56e-12 $X=11500 $Y=18000 $D=1
M1 GND A1 Y GND N L=4e-07 W=2e-06 AD=2.56e-12 AS=2.4e-12 $X=19500 $Y=18000 $D=1
M2 6 A0 VDD VDD P L=4e-07 W=5.2e-06 AD=3.12e-12 AS=5.98e-12 $X=11500 $Y=76000 $D=0
M3 Y A1 6 VDD P L=4e-07 W=5.2e-06 AD=5.62e-12 AS=3.12e-12 $X=16500 $Y=76000 $D=0
.ENDS
***************************************
.SUBCKT ICV_27 1
** N=2 EP=1 IP=4 FDC=80
X0 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
X1 1 2 ICV_19 $T=184000 0 0 0 $X=184000 $Y=0
.ENDS
***************************************
.SUBCKT ICV_28 1
** N=2 EP=1 IP=4 FDC=80
X0 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
X1 1 2 ICV_19 $T=0 0 1 180 $X=-244000 $Y=0
.ENDS
***************************************
.SUBCKT ao22 GND
** N=11 EP=1 IP=3 FDC=10
M0 10 B1 GND GND N L=4e-07 W=2e-06 AD=1.2e-12 AS=2.2e-12 $X=11500 $Y=26000 $D=1
M1 7 B0 10 GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=1.2e-12 $X=16500 $Y=26000 $D=1
M2 11 A0 7 GND N L=4e-07 W=2e-06 AD=1.2e-12 AS=2.4e-12 $X=24500 $Y=26000 $D=1
M3 GND A1 11 GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=1.2e-12 $X=29500 $Y=26000 $D=1
M4 Y 7 GND GND N L=4e-07 W=1e-06 AD=1.1e-12 AS=2.4e-12 $X=38000 $Y=31000 $D=1
M5 7 B1 8 VDD P L=4e-07 W=2.6e-06 AD=3.12e-12 AS=2.56e-12 $X=11500 $Y=76000 $D=0
M6 8 B0 7 VDD P L=4e-07 W=2.6e-06 AD=3.12e-12 AS=3.12e-12 $X=19500 $Y=76000 $D=0
M7 VDD A0 8 VDD P L=4e-07 W=2.6e-06 AD=3.12e-12 AS=3.12e-12 $X=27500 $Y=76000 $D=0
M8 8 A1 VDD VDD P L=4e-07 W=2.6e-06 AD=2.56e-12 AS=3.12e-12 $X=35500 $Y=76000 $D=0
M9 Y 7 VDD VDD P L=4e-07 W=1.8e-06 AD=1.58e-12 AS=1.58e-12 $X=51500 $Y=80000 $D=0
.ENDS
***************************************
.SUBCKT ICV_29 1
** N=2 EP=1 IP=4 FDC=76
X0 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
X1 1 2 ICV_16 $T=184000 0 0 0 $X=184000 $Y=0
.ENDS
***************************************
.SUBCKT aoi221 GND
** N=12 EP=1 IP=3 FDC=10
M0 Y C0 GND GND N L=4e-07 W=2e-06 AD=3.7e-12 AS=2.2e-12 $X=11500 $Y=26000 $D=1
M1 11 B0 Y GND N L=4e-07 W=3e-06 AD=1.8e-12 AS=3.7e-12 $X=20000 $Y=21000 $D=1
M2 GND B1 11 GND N L=4e-07 W=3e-06 AD=3.6e-12 AS=1.8e-12 $X=25000 $Y=21000 $D=1
M3 12 A1 GND GND N L=4e-07 W=3e-06 AD=1.8e-12 AS=3.6e-12 $X=33000 $Y=21000 $D=1
M4 Y A0 12 GND N L=4e-07 W=3e-06 AD=3.3e-12 AS=1.8e-12 $X=38000 $Y=21000 $D=1
M5 8 C0 Y VDD P L=4e-07 W=4.8e-06 AD=5.76e-12 AS=4.88e-12 $X=11500 $Y=73000 $D=0
M6 10 B0 8 VDD P L=4e-07 W=4.8e-06 AD=5.76e-12 AS=5.76e-12 $X=19500 $Y=73000 $D=0
M7 8 B1 10 VDD P L=4e-07 W=4.8e-06 AD=4.88e-12 AS=5.76e-12 $X=27500 $Y=73000 $D=0
M8 VDD A1 10 VDD P L=4e-07 W=4.8e-06 AD=5.76e-12 AS=4.88e-12 $X=44000 $Y=73000 $D=0
M9 10 A0 VDD VDD P L=4e-07 W=4.8e-06 AD=4.88e-12 AS=5.76e-12 $X=52000 $Y=73000 $D=0
.ENDS
***************************************
.SUBCKT oai21 GND VDD
** N=8 EP=2 IP=2 FDC=6
M0 7 B0 GND GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.2e-12 $X=11500 $Y=26000 $D=1
M1 Y A0 7 GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.4e-12 $X=19500 $Y=26000 $D=1
M2 7 A1 Y GND N L=4e-07 W=2e-06 AD=2.2e-12 AS=2.4e-12 $X=27500 $Y=26000 $D=1
M3 VDD B0 Y VDD P L=4e-07 W=2.4e-06 AD=5.76e-12 AS=2.44e-12 $X=11500 $Y=65000 $D=0
M4 8 A0 VDD VDD P L=4e-07 W=4.8e-06 AD=2.88e-12 AS=5.76e-12 $X=20000 $Y=65000 $D=0
M5 Y A1 8 VDD P L=4e-07 W=4.8e-06 AD=4.88e-12 AS=2.88e-12 $X=25000 $Y=65000 $D=0
.ENDS
***************************************
.SUBCKT nor03_2x GND
** N=8 EP=1 IP=0 FDC=6
M0 Y A0 GND GND N L=4e-07 W=2.2e-06 AD=2.64e-12 AS=2.68e-12 $X=11500 $Y=18000 $D=1
M1 GND A1 Y GND N L=4e-07 W=2.2e-06 AD=2.96e-12 AS=2.64e-12 $X=19500 $Y=18000 $D=1
M2 Y A2 GND GND N L=4e-07 W=2.2e-06 AD=2.32e-12 AS=2.96e-12 $X=27500 $Y=18000 $D=1
M3 7 A0 VDD VDD P L=4e-07 W=8e-06 AD=4.8e-12 AS=9.16e-12 $X=11500 $Y=62000 $D=0
M4 8 A1 7 VDD P L=4e-07 W=8e-06 AD=4.8e-12 AS=4.8e-12 $X=16500 $Y=62000 $D=0
M5 Y A2 8 VDD P L=4e-07 W=8e-06 AD=8.8e-12 AS=4.8e-12 $X=21500 $Y=62000 $D=0
.ENDS
***************************************
.SUBCKT inv04 GND
** N=4 EP=1 IP=1 FDC=4
M0 Y A GND GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.2e-12 $X=11500 $Y=26000 $D=1
M1 GND A Y GND N L=4e-07 W=2e-06 AD=2.2e-12 AS=2.4e-12 $X=19500 $Y=26000 $D=1
M2 Y A VDD VDD P L=4e-07 W=3.6e-06 AD=4.32e-12 AS=3.66e-12 $X=11500 $Y=71000 $D=0
M3 VDD A Y VDD P L=4e-07 W=3.6e-06 AD=3.66e-12 AS=4.32e-12 $X=19500 $Y=71000 $D=0
.ENDS
***************************************
.SUBCKT aoi21 GND
** N=8 EP=1 IP=2 FDC=6
M0 8 A1 GND GND N L=4e-07 W=2e-06 AD=1.2e-12 AS=2.2e-12 $X=11500 $Y=26000 $D=1
M1 Y A0 8 GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=1.2e-12 $X=16500 $Y=26000 $D=1
M2 GND B0 Y GND N L=4e-07 W=1e-06 AD=1.1e-12 AS=2.4e-12 $X=25000 $Y=31000 $D=1
M3 VDD A1 7 VDD P L=4e-07 W=2.6e-06 AD=3.12e-12 AS=2.56e-12 $X=11500 $Y=76000 $D=0
M4 7 A0 VDD VDD P L=4e-07 W=2.6e-06 AD=3.12e-12 AS=3.12e-12 $X=19500 $Y=76000 $D=0
M5 Y B0 7 VDD P L=4e-07 W=2.6e-06 AD=2.56e-12 AS=3.12e-12 $X=27500 $Y=76000 $D=0
.ENDS
***************************************
.SUBCKT ICV_30 1
** N=2 EP=1 IP=4 FDC=40
X0 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
X1 1 2 oai21 $T=184000 0 0 0 $X=184000 $Y=0
.ENDS
***************************************
.SUBCKT ICV_31 1
** N=2 EP=1 IP=4 FDC=42
X0 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
X1 1 2 nand04 $T=233000 0 1 180 $X=184000 $Y=0
.ENDS
***************************************
.SUBCKT ICV_32 1
** N=2 EP=1 IP=4 FDC=76
X0 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
X1 1 2 ICV_9 $T=184000 0 0 0 $X=184000 $Y=0
.ENDS
***************************************
.SUBCKT ICV_33 1
** N=2 EP=1 IP=4 FDC=40
X0 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
X1 1 2 oai21 $T=225000 0 1 180 $X=184000 $Y=0
.ENDS
***************************************
.SUBCKT ICV_34 1 2
** N=2 EP=2 IP=4 FDC=114
X0 1 2 ICV_4 $T=0 0 0 0 $X=0 $Y=0
X1 1 2 ICV_19 $T=368000 0 0 0 $X=368000 $Y=0
.ENDS
***************************************
.SUBCKT nor04 GND VDD
** N=10 EP=2 IP=3 FDC=8
M0 GND A3 Y GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.2e-12 $X=11500 $Y=21000 $D=1
M1 Y A2 GND GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.4e-12 $X=19500 $Y=21000 $D=1
M2 GND A1 Y GND N L=4e-07 W=2e-06 AD=2.4e-12 AS=2.4e-12 $X=27500 $Y=21000 $D=1
M3 Y A0 GND GND N L=4e-07 W=2e-06 AD=2.2e-12 AS=2.4e-12 $X=35500 $Y=21000 $D=1
M4 8 A3 Y VDD P L=4e-07 W=7.2e-06 AD=4.32e-12 AS=7.82e-12 $X=17500 $Y=69000 $D=0
M5 9 A2 8 VDD P L=4e-07 W=7.2e-06 AD=4.32e-12 AS=4.32e-12 $X=22500 $Y=69000 $D=0
M6 10 A1 9 VDD P L=4e-07 W=7.2e-06 AD=4.32e-12 AS=4.32e-12 $X=27500 $Y=69000 $D=0
M7 VDD A0 10 VDD P L=4e-07 W=7.2e-06 AD=7.82e-12 AS=4.32e-12 $X=32500 $Y=69000 $D=0
.ENDS
***************************************
.SUBCKT ICV_35 1
** N=2 EP=1 IP=4 FDC=36
X0 1 2 inv02 $T=0 0 1 180 $X=-25000 $Y=0
X1 1 2 dffr $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT or02 VDD GND
** N=7 EP=2 IP=2 FDC=6
M0 6 A1 GND GND N L=4e-07 W=1e-06 AD=1.2e-12 AS=1.1e-12 $X=11500 $Y=26000 $D=1
M1 GND A0 6 GND N L=4e-07 W=1e-06 AD=1.2e-12 AS=1.2e-12 $X=19500 $Y=26000 $D=1
M2 Y 6 GND GND N L=4e-07 W=1e-06 AD=1.1e-12 AS=1.2e-12 $X=27500 $Y=26000 $D=1
M3 7 A1 6 VDD P L=4e-07 W=2.6e-06 AD=1.56e-12 AS=2.56e-12 $X=11500 $Y=76000 $D=0
M4 VDD A0 7 VDD P L=4e-07 W=2.6e-06 AD=3.22e-12 AS=1.56e-12 $X=16500 $Y=76000 $D=0
M5 Y 6 VDD VDD P L=4e-07 W=1.8e-06 AD=1.58e-12 AS=3.22e-12 $X=25000 $Y=76000 $D=0
.ENDS
***************************************
.SUBCKT or03 GND VDD
** N=9 EP=2 IP=2 FDC=8
M0 GND 7 Y GND N L=4e-07 W=1e-06 AD=1.32e-12 AS=1.1e-12 $X=13500 $Y=26000 $D=1
M1 7 A2 GND GND N L=4e-07 W=1.2e-06 AD=1.44e-12 AS=1.32e-12 $X=21500 $Y=25000 $D=1
M2 GND A1 7 GND N L=4e-07 W=1.2e-06 AD=1.44e-12 AS=1.44e-12 $X=29500 $Y=25000 $D=1
M3 7 A0 GND GND N L=4e-07 W=1.2e-06 AD=1.22e-12 AS=1.44e-12 $X=37500 $Y=25000 $D=1
M4 VDD 7 Y VDD P L=4e-07 W=1.8e-06 AD=1.58e-12 AS=1.58e-12 $X=11500 $Y=80000 $D=0
M5 8 A2 7 VDD P L=4e-07 W=5.4e-06 AD=3.24e-12 AS=5.74e-12 $X=27500 $Y=73000 $D=0
M6 9 A1 8 VDD P L=4e-07 W=5.4e-06 AD=3.24e-12 AS=3.24e-12 $X=32500 $Y=73000 $D=0
M7 VDD A0 9 VDD P L=4e-07 W=5.4e-06 AD=5.74e-12 AS=3.24e-12 $X=37500 $Y=73000 $D=0
.ENDS
***************************************
.SUBCKT ICV_36 1
** N=3 EP=1 IP=4 FDC=18
X0 1 2 oai22 $T=-1000 0 1 180 $X=-50000 $Y=0
X1 1 3 xnor2 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_37 1
** N=3 EP=1 IP=4 FDC=12
X0 1 2 inv01 $T=-1000 0 1 180 $X=-26000 $Y=0
X1 1 3 xnor2 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT nand03 GND
** N=8 EP=1 IP=2 FDC=6
M0 7 A0 Y GND N L=4e-07 W=3e-06 AD=1.8e-12 AS=3.3e-12 $X=14500 $Y=26500 $D=1
M1 8 A1 7 GND N L=4e-07 W=3e-06 AD=1.8e-12 AS=1.8e-12 $X=19500 $Y=26500 $D=1
M2 GND A2 8 GND N L=4e-07 W=3e-06 AD=3.3e-12 AS=1.8e-12 $X=24500 $Y=26500 $D=1
M3 Y A0 VDD VDD P L=4e-07 W=3e-06 AD=3.6e-12 AS=3.3e-12 $X=11500 $Y=74000 $D=0
M4 VDD A1 Y VDD P L=4e-07 W=3e-06 AD=3.6e-12 AS=3.6e-12 $X=19500 $Y=74000 $D=0
M5 Y A2 VDD VDD P L=4e-07 W=3e-06 AD=3.3e-12 AS=3.6e-12 $X=27500 $Y=74000 $D=0
.ENDS
***************************************
.SUBCKT ao32 GND
** N=13 EP=1 IP=3 FDC=12
M0 GND 9 Y GND N L=4e-07 W=1e-06 AD=3.5e-12 AS=1.1e-12 $X=11500 $Y=36000 $D=1
M1 11 A2 GND GND N L=4e-07 W=3e-06 AD=1.8e-12 AS=3.5e-12 $X=20000 $Y=26000 $D=1
M2 12 A1 11 GND N L=4e-07 W=3e-06 AD=1.8e-12 AS=1.8e-12 $X=25000 $Y=26000 $D=1
M3 9 A0 12 GND N L=4e-07 W=3e-06 AD=3.7e-12 AS=1.8e-12 $X=30000 $Y=26000 $D=1
M4 13 B0 9 GND N L=4e-07 W=2e-06 AD=1.2e-12 AS=3.7e-12 $X=38500 $Y=26000 $D=1
M5 GND B1 13 GND N L=4e-07 W=2e-06 AD=2.2e-12 AS=1.2e-12 $X=43500 $Y=26000 $D=1
M6 VDD 9 Y VDD P L=4e-07 W=1.8e-06 AD=3.22e-12 AS=1.58e-12 $X=11500 $Y=76000 $D=0
M7 10 A2 VDD VDD P L=4e-07 W=2.6e-06 AD=3.12e-12 AS=3.22e-12 $X=20000 $Y=76000 $D=0
M8 VDD A1 10 VDD P L=4e-07 W=2.6e-06 AD=3.12e-12 AS=3.12e-12 $X=28000 $Y=76000 $D=0
M9 10 A0 VDD VDD P L=4e-07 W=2.6e-06 AD=3.12e-12 AS=3.12e-12 $X=36000 $Y=76000 $D=0
M10 9 B0 10 VDD P L=4e-07 W=2.6e-06 AD=3.12e-12 AS=3.12e-12 $X=44000 $Y=76000 $D=0
M11 10 B1 9 VDD P L=4e-07 W=2.6e-06 AD=2.56e-12 AS=3.12e-12 $X=52000 $Y=76000 $D=0
.ENDS
***************************************
.SUBCKT nor02ii GND
** N=7 EP=1 IP=0 FDC=6
M0 Y A0 GND GND N L=4e-07 W=1e-06 AD=1.2e-12 AS=1.1e-12 $X=11500 $Y=36000 $D=1
M1 GND 6 Y GND N L=4e-07 W=1e-06 AD=1.2e-12 AS=1.2e-12 $X=19500 $Y=36000 $D=1
M2 6 A1 GND GND N L=4e-07 W=1e-06 AD=1.1e-12 AS=1.2e-12 $X=27500 $Y=36000 $D=1
M3 7 A0 Y VDD P L=4e-07 W=2.6e-06 AD=1.56e-12 AS=2.56e-12 $X=11500 $Y=65000 $D=0
M4 VDD 6 7 VDD P L=4e-07 W=2.6e-06 AD=3.22e-12 AS=1.56e-12 $X=16500 $Y=65000 $D=0
M5 6 A1 VDD VDD P L=4e-07 W=1.8e-06 AD=1.58e-12 AS=3.22e-12 $X=25000 $Y=65000 $D=0
.ENDS
***************************************
.SUBCKT nand02_2x GND
** N=6 EP=1 IP=0 FDC=4
M0 6 A1 GND GND N L=4e-07 W=4e-06 AD=2.4e-12 AS=4.76e-12 $X=11500 $Y=18000 $D=1
M1 Y A0 6 GND N L=4e-07 W=4e-06 AD=4.4e-12 AS=2.4e-12 $X=16500 $Y=18000 $D=1
M2 Y A1 VDD VDD P L=4e-07 W=4e-06 AD=4.8e-12 AS=4.76e-12 $X=11500 $Y=82000 $D=0
M3 VDD A0 Y VDD P L=4e-07 W=4e-06 AD=4.76e-12 AS=4.8e-12 $X=19500 $Y=82000 $D=0
.ENDS
***************************************
.SUBCKT ICV_38 1
** N=3 EP=1 IP=4 FDC=18
X0 2 1 aoi22 $T=-50000 0 0 0 $X=-50000 $Y=0
X1 1 3 xnor2 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_39 1
** N=3 EP=1 IP=4 FDC=20
X0 1 2 xnor2 $T=-1000 0 1 180 $X=-64000 $Y=0
X1 1 3 xnor2 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT ICV_40 1
** N=3 EP=1 IP=4 FDC=18
X0 1 2 oai22 $T=64000 0 0 0 $X=64000 $Y=0
X1 1 3 xnor2 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
.SUBCKT system
** N=5835 EP=0 IP=12311 FDC=122912
X0 25 24 tri01 $T=10400000 96000 0 0 $X=10400000 $Y=96000
X1 26 24 tri01 $T=10400000 792000 0 0 $X=10400000 $Y=792000
X2 27 24 tri01 $T=10488000 328000 0 0 $X=10488000 $Y=328000
X3 28 24 tri01 $T=10504000 96000 0 0 $X=10504000 $Y=96000
X4 29 24 tri01 $T=10544000 96000 0 0 $X=10544000 $Y=96000
X5 30 24 tri01 $T=10630500 328000 1 180 $X=10592000 $Y=328000
X6 31 24 tri01 $T=10712000 96000 0 0 $X=10712000 $Y=96000
X7 32 24 tri01 $T=10774500 1488000 1 180 $X=10736000 $Y=1488000
X8 33 24 tri01 $T=10752000 96000 0 0 $X=10752000 $Y=96000
X9 34 24 tri01 $T=10920000 96000 0 0 $X=10920000 $Y=96000
X10 35 24 tri01 $T=10992000 1024000 0 0 $X=10992000 $Y=1024000
X11 36 24 tri01 $T=11016000 328000 0 0 $X=11016000 $Y=328000
X12 37 24 tri01 $T=11016000 1256000 0 0 $X=11016000 $Y=1256000
X13 38 24 tri01 $T=11062500 96000 1 180 $X=11024000 $Y=96000
X14 39 24 tri01 $T=11032000 1024000 0 0 $X=11032000 $Y=1024000
X15 40 24 tri01 $T=11056000 1256000 0 0 $X=11056000 $Y=1256000
X16 41 24 tri01 $T=11158500 328000 1 180 $X=11120000 $Y=328000
X17 42 24 tri01 $T=11136000 1024000 0 0 $X=11136000 $Y=1024000
X18 43 24 tri01 $T=11152000 792000 0 0 $X=11152000 $Y=792000
X19 44 24 tri01 $T=11152000 1488000 0 0 $X=11152000 $Y=1488000
X20 45 24 tri01 $T=11160000 328000 0 0 $X=11160000 $Y=328000
X21 46 24 tri01 $T=11160000 1256000 0 0 $X=11160000 $Y=1256000
X22 47 24 tri01 $T=11230500 96000 1 180 $X=11192000 $Y=96000
X23 48 24 tri01 $T=11262500 560000 1 180 $X=11224000 $Y=560000
X24 49 24 tri01 $T=11270500 96000 1 180 $X=11232000 $Y=96000
X25 50 24 tri01 $T=11294500 792000 1 180 $X=11256000 $Y=792000
X26 51 24 tri01 $T=11264000 328000 0 0 $X=11264000 $Y=328000
X27 52 24 tri01 $T=11264000 560000 0 0 $X=11264000 $Y=560000
X28 53 24 tri01 $T=11302500 1256000 1 180 $X=11264000 $Y=1256000
X29 54 24 tri01 $T=11272000 96000 0 0 $X=11272000 $Y=96000
X30 55 24 tri01 $T=11296000 792000 0 0 $X=11296000 $Y=792000
X31 56 24 tri01 $T=11304000 560000 0 0 $X=11304000 $Y=560000
X32 57 24 tri01 $T=11304000 1024000 0 0 $X=11304000 $Y=1024000
X33 58 24 tri01 $T=11312000 96000 0 0 $X=11312000 $Y=96000
X34 59 24 tri01 $T=11336000 792000 0 0 $X=11336000 $Y=792000
X35 60 24 tri01 $T=11344000 560000 0 0 $X=11344000 $Y=560000
X36 61 24 tri01 $T=11368000 328000 0 0 $X=11368000 $Y=328000
X37 62 24 tri01 $T=11376000 792000 0 0 $X=11376000 $Y=792000
X38 63 24 tri01 $T=11416000 96000 0 0 $X=11416000 $Y=96000
X39 64 24 tri01 $T=11456000 96000 0 0 $X=11456000 $Y=96000
X40 65 24 tri01 $T=11480000 1488000 0 0 $X=11480000 $Y=1488000
X41 66 24 tri01 $T=11512000 560000 0 0 $X=11512000 $Y=560000
X42 67 24 tri01 $T=11598500 96000 1 180 $X=11560000 $Y=96000
X43 68 24 tri01 $T=11598500 1256000 1 180 $X=11560000 $Y=1256000
X44 69 24 tri01 $T=11600000 96000 0 0 $X=11600000 $Y=96000
X45 70 24 tri01 $T=11608000 792000 0 0 $X=11608000 $Y=792000
X46 71 24 tri01 $T=11654500 560000 1 180 $X=11616000 $Y=560000
X47 72 24 tri01 $T=11640000 96000 0 0 $X=11640000 $Y=96000
X48 73 24 tri01 $T=11702500 1256000 1 180 $X=11664000 $Y=1256000
X49 74 24 tri01 $T=11702500 1488000 1 180 $X=11664000 $Y=1488000
X50 75 24 tri01 $T=11742500 1256000 1 180 $X=11704000 $Y=1256000
X51 76 24 tri01 $T=11750500 792000 1 180 $X=11712000 $Y=792000
X52 77 24 tri01 $T=11744000 1256000 0 0 $X=11744000 $Y=1256000
X53 78 24 tri01 $T=11752000 792000 0 0 $X=11752000 $Y=792000
X54 79 24 tri01 $T=11792000 792000 0 0 $X=11792000 $Y=792000
X55 80 24 tri01 $T=11838500 560000 1 180 $X=11800000 $Y=560000
X56 81 24 tri01 $T=11808000 96000 0 0 $X=11808000 $Y=96000
X57 82 24 tri01 $T=11808000 1488000 0 0 $X=11808000 $Y=1488000
X58 83 24 tri01 $T=11816000 7056000 0 0 $X=11816000 $Y=7056000
X59 84 24 tri01 $T=11862500 328000 1 180 $X=11824000 $Y=328000
X60 85 24 tri01 $T=11864000 328000 0 0 $X=11864000 $Y=328000
X61 86 24 tri01 $T=11904000 328000 0 0 $X=11904000 $Y=328000
X62 87 24 tri01 $T=11904000 8680000 0 0 $X=11904000 $Y=8680000
X63 88 24 tri01 $T=11950500 96000 1 180 $X=11912000 $Y=96000
X64 89 24 tri01 $T=11950500 1488000 1 180 $X=11912000 $Y=1488000
X65 90 24 tri01 $T=11936000 560000 0 0 $X=11936000 $Y=560000
X66 91 24 tri01 $T=11944000 1256000 0 0 $X=11944000 $Y=1256000
X67 92 24 tri01 $T=11952000 96000 0 0 $X=11952000 $Y=96000
X68 93 24 tri01 $T=11960000 792000 0 0 $X=11960000 $Y=792000
X69 94 24 tri01 $T=11968000 7288000 0 0 $X=11968000 $Y=7288000
X70 95 24 tri01 $T=11984000 1488000 0 0 $X=11984000 $Y=1488000
X71 96 24 tri01 $T=11992000 7056000 0 0 $X=11992000 $Y=7056000
X72 97 24 tri01 $T=12008000 7288000 0 0 $X=12008000 $Y=7288000
X73 98 24 tri01 $T=12078500 560000 1 180 $X=12040000 $Y=560000
X74 99 24 tri01 $T=12094500 96000 1 180 $X=12056000 $Y=96000
X75 100 24 tri01 $T=12064000 792000 0 0 $X=12064000 $Y=792000
X76 101 24 tri01 $T=12072000 8680000 0 0 $X=12072000 $Y=8680000
X77 102 24 tri01 $T=12096000 96000 0 0 $X=12096000 $Y=96000
X78 103 24 tri01 $T=12134500 7056000 1 180 $X=12096000 $Y=7056000
X79 104 24 tri01 $T=12136000 96000 0 0 $X=12136000 $Y=96000
X80 105 24 tri01 $T=12136000 328000 0 0 $X=12136000 $Y=328000
X81 106 24 tri01 $T=12174500 7520000 1 180 $X=12136000 $Y=7520000
X82 107 24 tri01 $T=12144000 1024000 0 0 $X=12144000 $Y=1024000
X83 108 24 tri01 $T=12176000 96000 0 0 $X=12176000 $Y=96000
X84 109 24 tri01 $T=12176000 1256000 0 0 $X=12176000 $Y=1256000
X85 110 24 tri01 $T=12176000 7520000 0 0 $X=12176000 $Y=7520000
X86 111 24 tri01 $T=12214500 8912000 1 180 $X=12176000 $Y=8912000
X87 112 24 tri01 $T=12200000 792000 0 0 $X=12200000 $Y=792000
X88 113 24 tri01 $T=12240000 7288000 0 0 $X=12240000 $Y=7288000
X89 114 24 tri01 $T=12286500 1024000 1 180 $X=12248000 $Y=1024000
X90 115 24 tri01 $T=12318500 1256000 1 180 $X=12280000 $Y=1256000
X91 116 24 tri01 $T=12318500 1488000 1 180 $X=12280000 $Y=1488000
X92 117 24 tri01 $T=12318500 7520000 1 180 $X=12280000 $Y=7520000
X93 118 24 tri01 $T=12342500 792000 1 180 $X=12304000 $Y=792000
X94 119 24 tri01 $T=12320000 1488000 0 0 $X=12320000 $Y=1488000
X95 120 24 tri01 $T=12382500 96000 1 180 $X=12344000 $Y=96000
X96 121 24 tri01 $T=12344000 328000 0 0 $X=12344000 $Y=328000
X97 122 24 tri01 $T=12344000 792000 0 0 $X=12344000 $Y=792000
X98 123 24 tri01 $T=12382500 7288000 1 180 $X=12344000 $Y=7288000
X99 124 24 tri01 $T=12344000 8912000 0 0 $X=12344000 $Y=8912000
X100 125 24 tri01 $T=12414500 1720000 1 180 $X=12376000 $Y=1720000
X101 126 24 tri01 $T=12384000 7288000 0 0 $X=12384000 $Y=7288000
X102 127 24 tri01 $T=12454500 1024000 1 180 $X=12416000 $Y=1024000
X103 128 24 tri01 $T=12486500 96000 1 180 $X=12448000 $Y=96000
X104 129 24 tri01 $T=12486500 328000 1 180 $X=12448000 $Y=328000
X105 130 24 tri01 $T=12486500 792000 1 180 $X=12448000 $Y=792000
X106 131 24 tri01 $T=12486500 1256000 1 180 $X=12448000 $Y=1256000
X107 132 24 tri01 $T=12448000 1720000 0 0 $X=12448000 $Y=1720000
X108 133 24 tri01 $T=12486500 6824000 1 180 $X=12448000 $Y=6824000
X109 134 24 tri01 $T=12486500 7520000 1 180 $X=12448000 $Y=7520000
X110 135 24 tri01 $T=12486500 8912000 1 180 $X=12448000 $Y=8912000
X111 136 24 tri01 $T=12526500 96000 1 180 $X=12488000 $Y=96000
X112 137 24 tri01 $T=12526500 328000 1 180 $X=12488000 $Y=328000
X113 138 24 tri01 $T=12526500 560000 1 180 $X=12488000 $Y=560000
X114 139 24 tri01 $T=12526500 792000 1 180 $X=12488000 $Y=792000
X115 140 24 tri01 $T=12526500 1024000 1 180 $X=12488000 $Y=1024000
X116 141 24 tri01 $T=12526500 1256000 1 180 $X=12488000 $Y=1256000
X117 142 24 tri01 $T=12526500 1488000 1 180 $X=12488000 $Y=1488000
X118 143 24 tri01 $T=12526500 6824000 1 180 $X=12488000 $Y=6824000
X119 144 24 tri01 $T=12526500 7056000 1 180 $X=12488000 $Y=7056000
X120 145 24 tri01 $T=12526500 7288000 1 180 $X=12488000 $Y=7288000
X121 146 24 tri01 $T=12526500 7520000 1 180 $X=12488000 $Y=7520000
X122 147 24 tri01 $T=12526500 8680000 1 180 $X=12488000 $Y=8680000
X123 148 24 tri01 $T=12526500 8912000 1 180 $X=12488000 $Y=8912000
X124 24 nand02 $T=488000 8448000 0 0 $X=488000 $Y=8448000
X125 24 nand02 $T=488000 8680000 0 0 $X=488000 $Y=8680000
X126 24 nand02 $T=560000 8448000 0 0 $X=560000 $Y=8448000
X127 24 nand02 $T=600000 8448000 0 0 $X=600000 $Y=8448000
X128 24 nand02 $T=656000 8680000 0 0 $X=656000 $Y=8680000
X129 24 nand02 $T=672000 8448000 0 0 $X=672000 $Y=8448000
X130 24 nand02 $T=712000 8448000 0 0 $X=712000 $Y=8448000
X131 24 nand02 $T=736000 8680000 0 0 $X=736000 $Y=8680000
X132 24 nand02 $T=752000 8448000 0 0 $X=752000 $Y=8448000
X133 24 nand02 $T=760000 8912000 0 0 $X=760000 $Y=8912000
X134 24 nand02 $T=792000 8448000 0 0 $X=792000 $Y=8448000
X135 24 nand02 $T=808000 8680000 0 0 $X=808000 $Y=8680000
X136 24 nand02 $T=896000 8680000 0 0 $X=896000 $Y=8680000
X137 24 nand02 $T=896000 8912000 0 0 $X=896000 $Y=8912000
X138 24 nand02 $T=1433000 9840000 1 180 $X=1400000 $Y=9840000
X139 24 nand02 $T=1408000 10072000 0 0 $X=1408000 $Y=10072000
X140 24 nand02 $T=1481000 10072000 1 180 $X=1448000 $Y=10072000
X141 24 nand02 $T=1521000 10072000 1 180 $X=1488000 $Y=10072000
X142 24 nand02 $T=1576000 9840000 0 0 $X=1576000 $Y=9840000
X143 24 nand02 $T=1624000 10072000 0 0 $X=1624000 $Y=10072000
X144 24 nand02 $T=1704000 10072000 0 0 $X=1704000 $Y=10072000
X145 24 nand02 $T=1912000 10072000 0 0 $X=1912000 $Y=10072000
X146 24 nand02 $T=1961000 2880000 1 180 $X=1928000 $Y=2880000
X147 24 nand02 $T=2016000 10072000 0 0 $X=2016000 $Y=10072000
X148 24 nand02 $T=2160000 10072000 0 0 $X=2160000 $Y=10072000
X149 24 nand02 $T=2200000 10072000 0 0 $X=2200000 $Y=10072000
X150 24 nand02 $T=2304000 10072000 0 0 $X=2304000 $Y=10072000
X151 24 nand02 $T=2344000 10072000 0 0 $X=2344000 $Y=10072000
X152 24 nand02 $T=2384000 9840000 0 0 $X=2384000 $Y=9840000
X153 24 nand02 $T=2384000 10072000 0 0 $X=2384000 $Y=10072000
X154 24 nand02 $T=2424000 10072000 0 0 $X=2424000 $Y=10072000
X155 24 nand02 $T=2464000 10072000 0 0 $X=2464000 $Y=10072000
X156 24 nand02 $T=2569000 3112000 1 180 $X=2536000 $Y=3112000
X157 24 nand02 $T=2656000 2880000 0 0 $X=2656000 $Y=2880000
X158 24 nand02 $T=10440000 792000 0 0 $X=10440000 $Y=792000
X159 24 nand02 $T=10592000 1488000 0 0 $X=10592000 $Y=1488000
X160 24 nand02 $T=11176000 1024000 0 0 $X=11176000 $Y=1024000
X161 24 nand02 $T=11520000 1488000 0 0 $X=11520000 $Y=1488000
X162 24 nand02 $T=11656000 560000 0 0 $X=11656000 $Y=560000
X163 24 nand02 $T=11737000 1488000 1 180 $X=11704000 $Y=1488000
X164 24 nand02 $T=11817000 328000 1 180 $X=11784000 $Y=328000
X165 24 nand02 $T=11784000 1256000 0 0 $X=11784000 $Y=1256000
X166 24 nand02 $T=11856000 7288000 0 0 $X=11856000 $Y=7288000
X167 24 nand02 $T=11929000 6824000 1 180 $X=11896000 $Y=6824000
X168 24 nand02 $T=11984000 1024000 0 0 $X=11984000 $Y=1024000
X169 24 nand02 $T=12024000 1488000 0 0 $X=12024000 $Y=1488000
X170 24 nand02 $T=12137000 792000 1 180 $X=12104000 $Y=792000
X171 24 nand02 $T=12241000 1488000 1 180 $X=12208000 $Y=1488000
X172 24 nand02 $T=12304000 328000 0 0 $X=12304000 $Y=328000
X173 24 nand02 $T=12488000 1720000 0 0 $X=12488000 $Y=1720000
X174 24 149 oai22 $T=400000 4040000 0 0 $X=400000 $Y=4040000
X175 24 150 oai22 $T=505000 4040000 1 180 $X=456000 $Y=4040000
X176 24 151 oai22 $T=632000 4040000 0 0 $X=632000 $Y=4040000
X177 24 152 oai22 $T=697000 2416000 1 180 $X=648000 $Y=2416000
X178 24 153 oai22 $T=848000 3808000 0 0 $X=848000 $Y=3808000
X179 24 154 oai22 $T=905000 2880000 1 180 $X=856000 $Y=2880000
X180 24 155 oai22 $T=1048000 96000 0 0 $X=1048000 $Y=96000
X181 24 156 oai22 $T=1201000 2648000 1 180 $X=1152000 $Y=2648000
X182 24 157 oai22 $T=1416000 792000 0 0 $X=1416000 $Y=792000
X183 24 158 oai22 $T=1881000 2648000 1 180 $X=1832000 $Y=2648000
X184 24 159 oai22 $T=1880000 328000 0 0 $X=1880000 $Y=328000
X185 24 160 oai22 $T=1952000 2184000 0 0 $X=1952000 $Y=2184000
X186 24 161 oai22 $T=2104000 792000 0 0 $X=2104000 $Y=792000
X187 24 162 oai22 $T=2152000 560000 0 0 $X=2152000 $Y=560000
X188 24 163 oai22 $T=2401000 1720000 1 180 $X=2352000 $Y=1720000
X189 24 164 oai22 $T=2656000 2416000 0 0 $X=2656000 $Y=2416000
X190 24 165 oai22 $T=2904000 2880000 0 0 $X=2904000 $Y=2880000
X191 24 166 oai22 $T=2944000 1488000 0 0 $X=2944000 $Y=1488000
X192 24 167 oai22 $T=3065000 328000 1 180 $X=3016000 $Y=328000
X193 24 168 oai22 $T=4080000 328000 0 0 $X=4080000 $Y=328000
X194 24 169 oai22 $T=10561000 792000 1 180 $X=10512000 $Y=792000
X195 24 170 oai22 $T=10776000 1024000 0 0 $X=10776000 $Y=1024000
X196 24 171 oai22 $T=11216000 1024000 0 0 $X=11216000 $Y=1024000
X197 24 172 oai22 $T=11560000 6592000 0 0 $X=11560000 $Y=6592000
X198 24 173 oai22 $T=11728000 328000 0 0 $X=11728000 $Y=328000
X199 24 174 oai22 $T=11824000 1256000 0 0 $X=11824000 $Y=1256000
X200 24 175 oai22 $T=12024000 1024000 0 0 $X=12024000 $Y=1024000
X201 24 176 oai22 $T=12193000 792000 1 180 $X=12144000 $Y=792000
X202 24 177 oai22 $T=12336000 560000 0 0 $X=12336000 $Y=560000
X203 24 178 oai22 $T=12472000 1952000 0 0 $X=12472000 $Y=1952000
X204 24 179 inv02 $T=369000 2648000 1 180 $X=344000 $Y=2648000
X205 24 180 inv02 $T=369000 3112000 1 180 $X=344000 $Y=3112000
X206 24 181 inv02 $T=401000 3112000 1 180 $X=376000 $Y=3112000
X207 24 182 inv02 $T=465000 10768000 1 180 $X=440000 $Y=10768000
X208 24 183 inv02 $T=440000 12392000 0 0 $X=440000 $Y=12392000
X209 24 184 inv02 $T=440000 12624000 0 0 $X=440000 $Y=12624000
X210 24 185 inv02 $T=472000 10768000 0 0 $X=472000 $Y=10768000
X211 24 186 inv02 $T=472000 12624000 0 0 $X=472000 $Y=12624000
X212 24 187 inv02 $T=480000 12160000 0 0 $X=480000 $Y=12160000
X213 24 188 inv02 $T=504000 7520000 0 0 $X=504000 $Y=7520000
X214 24 189 inv02 $T=528000 8448000 0 0 $X=528000 $Y=8448000
X215 24 190 inv02 $T=536000 1720000 0 0 $X=536000 $Y=1720000
X216 24 191 inv02 $T=577000 10072000 1 180 $X=552000 $Y=10072000
X217 24 192 inv02 $T=577000 12160000 1 180 $X=552000 $Y=12160000
X218 24 193 inv02 $T=585000 10768000 1 180 $X=560000 $Y=10768000
X219 24 194 inv02 $T=584000 10072000 0 0 $X=584000 $Y=10072000
X220 24 195 inv02 $T=584000 12160000 0 0 $X=584000 $Y=12160000
X221 24 196 inv02 $T=641000 12160000 1 180 $X=616000 $Y=12160000
X222 24 197 inv02 $T=624000 8680000 0 0 $X=624000 $Y=8680000
X223 24 198 inv02 $T=640000 8448000 0 0 $X=640000 $Y=8448000
X224 24 199 inv02 $T=648000 12160000 0 0 $X=648000 $Y=12160000
X225 24 200 inv02 $T=672000 328000 0 0 $X=672000 $Y=328000
X226 24 201 inv02 $T=672000 10768000 0 0 $X=672000 $Y=10768000
X227 24 202 inv02 $T=713000 7984000 1 180 $X=688000 $Y=7984000
X228 24 203 inv02 $T=721000 3808000 1 180 $X=696000 $Y=3808000
X229 24 204 inv02 $T=729000 9376000 1 180 $X=704000 $Y=9376000
X230 24 205 inv02 $T=712000 4272000 0 0 $X=712000 $Y=4272000
X231 24 206 inv02 $T=712000 7056000 0 0 $X=712000 $Y=7056000
X232 24 207 inv02 $T=712000 11928000 0 0 $X=712000 $Y=11928000
X233 24 208 inv02 $T=753000 1488000 1 180 $X=728000 $Y=1488000
X234 24 209 inv02 $T=761000 9376000 1 180 $X=736000 $Y=9376000
X235 24 210 inv02 $T=744000 4272000 0 0 $X=744000 $Y=4272000
X236 24 211 inv02 $T=785000 1488000 1 180 $X=760000 $Y=1488000
X237 24 212 inv02 $T=760000 11000000 0 0 $X=760000 $Y=11000000
X238 24 213 inv02 $T=801000 8680000 1 180 $X=776000 $Y=8680000
X239 24 214 inv02 $T=817000 1488000 1 180 $X=792000 $Y=1488000
X240 24 215 inv02 $T=792000 12160000 0 0 $X=792000 $Y=12160000
X241 24 216 inv02 $T=825000 6360000 1 180 $X=800000 $Y=6360000
X242 24 217 inv02 $T=825000 7520000 1 180 $X=800000 $Y=7520000
X243 24 218 inv02 $T=816000 1024000 0 0 $X=816000 $Y=1024000
X244 24 219 inv02 $T=849000 1488000 1 180 $X=824000 $Y=1488000
X245 24 220 inv02 $T=849000 5432000 1 180 $X=824000 $Y=5432000
X246 24 221 inv02 $T=849000 7984000 1 180 $X=824000 $Y=7984000
X247 24 222 inv02 $T=857000 6360000 1 180 $X=832000 $Y=6360000
X248 24 223 inv02 $T=832000 8448000 0 0 $X=832000 $Y=8448000
X249 24 224 inv02 $T=832000 10072000 0 0 $X=832000 $Y=10072000
X250 24 225 inv02 $T=848000 9376000 0 0 $X=848000 $Y=9376000
X251 24 226 inv02 $T=856000 7752000 0 0 $X=856000 $Y=7752000
X252 24 227 inv02 $T=880000 9144000 0 0 $X=880000 $Y=9144000
X253 24 228 inv02 $T=896000 3344000 0 0 $X=896000 $Y=3344000
X254 24 229 inv02 $T=896000 6824000 0 0 $X=896000 $Y=6824000
X255 24 230 inv02 $T=928000 6824000 0 0 $X=928000 $Y=6824000
X256 24 231 inv02 $T=936000 8680000 0 0 $X=936000 $Y=8680000
X257 24 232 inv02 $T=952000 9144000 0 0 $X=952000 $Y=9144000
X258 24 233 inv02 $T=968000 8680000 0 0 $X=968000 $Y=8680000
X259 24 234 inv02 $T=1040000 8680000 0 0 $X=1040000 $Y=8680000
X260 24 235 inv02 $T=1081000 4272000 1 180 $X=1056000 $Y=4272000
X261 24 236 inv02 $T=1105000 7520000 1 180 $X=1080000 $Y=7520000
X262 24 237 inv02 $T=1121000 1720000 1 180 $X=1096000 $Y=1720000
X263 24 238 inv02 $T=1161000 1256000 1 180 $X=1136000 $Y=1256000
X264 24 239 inv02 $T=1161000 8448000 1 180 $X=1136000 $Y=8448000
X265 24 240 inv02 $T=1193000 1256000 1 180 $X=1168000 $Y=1256000
X266 24 241 inv02 $T=1192000 10768000 0 0 $X=1192000 $Y=10768000
X267 24 242 inv02 $T=1200000 792000 0 0 $X=1200000 $Y=792000
X268 24 243 inv02 $T=1200000 1256000 0 0 $X=1200000 $Y=1256000
X269 24 244 inv02 $T=1200000 4040000 0 0 $X=1200000 $Y=4040000
X270 24 245 inv02 $T=1225000 5200000 1 180 $X=1200000 $Y=5200000
X271 24 246 inv02 $T=1200000 6128000 0 0 $X=1200000 $Y=6128000
X272 24 247 inv02 $T=1241000 10536000 1 180 $X=1216000 $Y=10536000
X273 24 248 inv02 $T=1257000 5200000 1 180 $X=1232000 $Y=5200000
X274 24 249 inv02 $T=1248000 3112000 0 0 $X=1248000 $Y=3112000
X275 24 250 inv02 $T=1289000 560000 1 180 $X=1264000 $Y=560000
X276 24 251 inv02 $T=1264000 2416000 0 0 $X=1264000 $Y=2416000
X277 24 252 inv02 $T=1296000 560000 0 0 $X=1296000 $Y=560000
X278 24 253 inv02 $T=1296000 2416000 0 0 $X=1296000 $Y=2416000
X279 24 254 inv02 $T=1296000 5432000 0 0 $X=1296000 $Y=5432000
X280 24 255 inv02 $T=1321000 10072000 1 180 $X=1296000 $Y=10072000
X281 24 256 inv02 $T=1345000 5896000 1 180 $X=1320000 $Y=5896000
X282 24 257 inv02 $T=1353000 2880000 1 180 $X=1328000 $Y=2880000
X283 24 258 inv02 $T=1344000 11232000 0 0 $X=1344000 $Y=11232000
X284 24 259 inv02 $T=1377000 13088000 1 180 $X=1352000 $Y=13088000
X285 24 260 inv02 $T=1360000 1024000 0 0 $X=1360000 $Y=1024000
X286 24 261 inv02 $T=1368000 2648000 0 0 $X=1368000 $Y=2648000
X287 24 262 inv02 $T=1368000 7056000 0 0 $X=1368000 $Y=7056000
X288 24 263 inv02 $T=1392000 9608000 0 0 $X=1392000 $Y=9608000
X289 24 264 inv02 $T=1400000 7056000 0 0 $X=1400000 $Y=7056000
X290 24 265 inv02 $T=1424000 9608000 0 0 $X=1424000 $Y=9608000
X291 24 266 inv02 $T=1456000 7288000 0 0 $X=1456000 $Y=7288000
X292 24 267 inv02 $T=1521000 1488000 1 180 $X=1496000 $Y=1488000
X293 24 268 inv02 $T=1528000 1488000 0 0 $X=1528000 $Y=1488000
X294 24 269 inv02 $T=1561000 3112000 1 180 $X=1536000 $Y=3112000
X295 24 270 inv02 $T=1569000 2648000 1 180 $X=1544000 $Y=2648000
X296 24 271 inv02 $T=1577000 2416000 1 180 $X=1552000 $Y=2416000
X297 24 272 inv02 $T=1552000 8448000 0 0 $X=1552000 $Y=8448000
X298 24 273 inv02 $T=1585000 1488000 1 180 $X=1560000 $Y=1488000
X299 24 274 inv02 $T=1568000 3576000 0 0 $X=1568000 $Y=3576000
X300 24 275 inv02 $T=1576000 5432000 0 0 $X=1576000 $Y=5432000
X301 24 276 inv02 $T=1609000 2416000 1 180 $X=1584000 $Y=2416000
X302 24 277 inv02 $T=1617000 1488000 1 180 $X=1592000 $Y=1488000
X303 24 278 inv02 $T=1641000 2416000 1 180 $X=1616000 $Y=2416000
X304 24 279 inv02 $T=1616000 11928000 0 0 $X=1616000 $Y=11928000
X305 24 280 inv02 $T=1649000 1488000 1 180 $X=1624000 $Y=1488000
X306 24 281 inv02 $T=1648000 2416000 0 0 $X=1648000 $Y=2416000
X307 24 282 inv02 $T=1673000 10536000 1 180 $X=1648000 $Y=10536000
X308 24 283 inv02 $T=1648000 11928000 0 0 $X=1648000 $Y=11928000
X309 24 284 inv02 $T=1656000 1488000 0 0 $X=1656000 $Y=1488000
X310 24 285 inv02 $T=1697000 10304000 1 180 $X=1672000 $Y=10304000
X311 24 286 inv02 $T=1680000 1720000 0 0 $X=1680000 $Y=1720000
X312 24 287 inv02 $T=1680000 1952000 0 0 $X=1680000 $Y=1952000
X313 24 288 inv02 $T=1680000 10536000 0 0 $X=1680000 $Y=10536000
X314 24 289 inv02 $T=1688000 1488000 0 0 $X=1688000 $Y=1488000
X315 24 290 inv02 $T=1713000 3112000 1 180 $X=1688000 $Y=3112000
X316 24 291 inv02 $T=1737000 1952000 1 180 $X=1712000 $Y=1952000
X317 24 292 inv02 $T=1720000 2184000 0 0 $X=1720000 $Y=2184000
X318 24 293 inv02 $T=1896000 4272000 0 0 $X=1896000 $Y=4272000
X319 24 294 inv02 $T=1921000 8680000 1 180 $X=1896000 $Y=8680000
X320 24 295 inv02 $T=1953000 4272000 1 180 $X=1928000 $Y=4272000
X321 24 296 inv02 $T=1952000 10072000 0 0 $X=1952000 $Y=10072000
X322 24 297 inv02 $T=1984000 7288000 0 0 $X=1984000 $Y=7288000
X323 24 298 inv02 $T=2009000 10072000 1 180 $X=1984000 $Y=10072000
X324 24 299 inv02 $T=1984000 10304000 0 0 $X=1984000 $Y=10304000
X325 24 300 inv02 $T=2017000 2648000 1 180 $X=1992000 $Y=2648000
X326 24 301 inv02 $T=1992000 7520000 0 0 $X=1992000 $Y=7520000
X327 24 302 inv02 $T=2016000 10304000 0 0 $X=2016000 $Y=10304000
X328 24 303 inv02 $T=2049000 11232000 1 180 $X=2024000 $Y=11232000
X329 24 304 inv02 $T=2048000 2184000 0 0 $X=2048000 $Y=2184000
X330 24 305 inv02 $T=2056000 10072000 0 0 $X=2056000 $Y=10072000
X331 24 306 inv02 $T=2113000 3112000 1 180 $X=2088000 $Y=3112000
X332 24 307 inv02 $T=2113000 9376000 1 180 $X=2088000 $Y=9376000
X333 24 308 inv02 $T=2145000 3112000 1 180 $X=2120000 $Y=3112000
X334 24 309 inv02 $T=2128000 10072000 0 0 $X=2128000 $Y=10072000
X335 24 310 inv02 $T=2153000 11000000 1 180 $X=2128000 $Y=11000000
X336 24 311 inv02 $T=2136000 12624000 0 0 $X=2136000 $Y=12624000
X337 24 312 inv02 $T=2144000 10304000 0 0 $X=2144000 $Y=10304000
X338 24 313 inv02 $T=2169000 11696000 1 180 $X=2144000 $Y=11696000
X339 24 314 inv02 $T=2177000 3112000 1 180 $X=2152000 $Y=3112000
X340 24 315 inv02 $T=2160000 11000000 0 0 $X=2160000 $Y=11000000
X341 24 316 inv02 $T=2193000 12624000 1 180 $X=2168000 $Y=12624000
X342 24 317 inv02 $T=2201000 10304000 1 180 $X=2176000 $Y=10304000
X343 24 318 inv02 $T=2200000 12624000 0 0 $X=2200000 $Y=12624000
X344 24 319 inv02 $T=2257000 3112000 1 180 $X=2232000 $Y=3112000
X345 24 320 inv02 $T=2257000 6824000 1 180 $X=2232000 $Y=6824000
X346 24 321 inv02 $T=2257000 11696000 1 180 $X=2232000 $Y=11696000
X347 24 322 inv02 $T=2257000 12624000 1 180 $X=2232000 $Y=12624000
X348 24 323 inv02 $T=2240000 10072000 0 0 $X=2240000 $Y=10072000
X349 24 324 inv02 $T=2289000 12624000 1 180 $X=2264000 $Y=12624000
X350 24 325 inv02 $T=2272000 10072000 0 0 $X=2272000 $Y=10072000
X351 24 326 inv02 $T=2305000 9144000 1 180 $X=2280000 $Y=9144000
X352 24 327 inv02 $T=2321000 3112000 1 180 $X=2296000 $Y=3112000
X353 24 328 inv02 $T=2321000 12624000 1 180 $X=2296000 $Y=12624000
X354 24 329 inv02 $T=2361000 2880000 1 180 $X=2336000 $Y=2880000
X355 24 330 inv02 $T=2361000 11928000 1 180 $X=2336000 $Y=11928000
X356 24 331 inv02 $T=2352000 2184000 0 0 $X=2352000 $Y=2184000
X357 24 332 inv02 $T=2352000 9840000 0 0 $X=2352000 $Y=9840000
X358 24 333 inv02 $T=2360000 2416000 0 0 $X=2360000 $Y=2416000
X359 24 334 inv02 $T=2385000 10536000 1 180 $X=2360000 $Y=10536000
X360 24 335 inv02 $T=2393000 11928000 1 180 $X=2368000 $Y=11928000
X361 24 336 inv02 $T=2409000 11232000 1 180 $X=2384000 $Y=11232000
X362 24 337 inv02 $T=2392000 2416000 0 0 $X=2392000 $Y=2416000
X363 24 338 inv02 $T=2432000 2184000 0 0 $X=2432000 $Y=2184000
X364 24 339 inv02 $T=2456000 3112000 0 0 $X=2456000 $Y=3112000
X365 24 340 inv02 $T=2497000 2880000 1 180 $X=2472000 $Y=2880000
X366 24 341 inv02 $T=2505000 12856000 1 180 $X=2480000 $Y=12856000
X367 24 342 inv02 $T=2488000 4272000 0 0 $X=2488000 $Y=4272000
X368 24 343 inv02 $T=2521000 10768000 1 180 $X=2496000 $Y=10768000
X369 24 344 inv02 $T=2537000 8448000 1 180 $X=2512000 $Y=8448000
X370 24 345 inv02 $T=2512000 11696000 0 0 $X=2512000 $Y=11696000
X371 24 346 inv02 $T=2537000 12856000 1 180 $X=2512000 $Y=12856000
X372 24 347 inv02 $T=2544000 7520000 0 0 $X=2544000 $Y=7520000
X373 24 348 inv02 $T=2544000 8448000 0 0 $X=2544000 $Y=8448000
X374 24 349 inv02 $T=2609000 2648000 1 180 $X=2584000 $Y=2648000
X375 24 350 inv02 $T=2625000 11696000 1 180 $X=2600000 $Y=11696000
X376 24 351 inv02 $T=2648000 12856000 0 0 $X=2648000 $Y=12856000
X377 24 352 inv02 $T=2689000 12624000 1 180 $X=2664000 $Y=12624000
X378 24 353 inv02 $T=2688000 11696000 0 0 $X=2688000 $Y=11696000
X379 24 354 inv02 $T=2752000 6360000 0 0 $X=2752000 $Y=6360000
X380 24 355 inv02 $T=2785000 10072000 1 180 $X=2760000 $Y=10072000
X381 24 356 inv02 $T=2793000 9376000 1 180 $X=2768000 $Y=9376000
X382 24 357 inv02 $T=2849000 328000 1 180 $X=2824000 $Y=328000
X383 24 358 inv02 $T=2857000 10768000 1 180 $X=2832000 $Y=10768000
X384 24 359 inv02 $T=2897000 11464000 1 180 $X=2872000 $Y=11464000
X385 24 360 inv02 $T=2945000 9840000 1 180 $X=2920000 $Y=9840000
X386 24 361 inv02 $T=2936000 11000000 0 0 $X=2936000 $Y=11000000
X387 24 362 inv02 $T=2977000 9840000 1 180 $X=2952000 $Y=9840000
X388 24 363 inv02 $T=2985000 9144000 1 180 $X=2960000 $Y=9144000
X389 24 364 inv02 $T=3001000 6824000 1 180 $X=2976000 $Y=6824000
X390 24 365 inv02 $T=2984000 11464000 0 0 $X=2984000 $Y=11464000
X391 24 366 inv02 $T=3017000 9144000 1 180 $X=2992000 $Y=9144000
X392 24 367 inv02 $T=3049000 11000000 1 180 $X=3024000 $Y=11000000
X393 24 368 inv02 $T=3065000 10072000 1 180 $X=3040000 $Y=10072000
X394 24 369 inv02 $T=3097000 7520000 1 180 $X=3072000 $Y=7520000
X395 24 370 inv02 $T=3097000 10072000 1 180 $X=3072000 $Y=10072000
X396 24 371 inv02 $T=3121000 2648000 1 180 $X=3096000 $Y=2648000
X397 24 372 inv02 $T=3096000 6360000 0 0 $X=3096000 $Y=6360000
X398 24 373 inv02 $T=3137000 4968000 1 180 $X=3112000 $Y=4968000
X399 24 374 inv02 $T=3120000 792000 0 0 $X=3120000 $Y=792000
X400 24 375 inv02 $T=3177000 8216000 1 180 $X=3152000 $Y=8216000
X401 24 376 inv02 $T=3160000 1488000 0 0 $X=3160000 $Y=1488000
X402 24 377 inv02 $T=3168000 7288000 0 0 $X=3168000 $Y=7288000
X403 24 378 inv02 $T=3209000 8448000 1 180 $X=3184000 $Y=8448000
X404 24 379 inv02 $T=3225000 7288000 1 180 $X=3200000 $Y=7288000
X405 24 380 inv02 $T=3232000 7288000 0 0 $X=3232000 $Y=7288000
X406 24 381 inv02 $T=3257000 10768000 1 180 $X=3232000 $Y=10768000
X407 24 382 inv02 $T=3256000 6824000 0 0 $X=3256000 $Y=6824000
X408 24 383 inv02 $T=3289000 10768000 1 180 $X=3264000 $Y=10768000
X409 24 384 inv02 $T=3288000 9840000 0 0 $X=3288000 $Y=9840000
X410 24 385 inv02 $T=3377000 10768000 1 180 $X=3352000 $Y=10768000
X411 24 386 inv02 $T=3384000 10768000 0 0 $X=3384000 $Y=10768000
X412 24 387 inv02 $T=3392000 5200000 0 0 $X=3392000 $Y=5200000
X413 24 388 inv02 $T=3416000 10768000 0 0 $X=3416000 $Y=10768000
X414 24 389 inv02 $T=3424000 10072000 0 0 $X=3424000 $Y=10072000
X415 24 390 inv02 $T=3473000 6592000 1 180 $X=3448000 $Y=6592000
X416 24 391 inv02 $T=3472000 8680000 0 0 $X=3472000 $Y=8680000
X417 24 392 inv02 $T=3593000 6824000 1 180 $X=3568000 $Y=6824000
X418 24 393 inv02 $T=3600000 6824000 0 0 $X=3600000 $Y=6824000
X419 24 394 inv02 $T=3673000 7056000 1 180 $X=3648000 $Y=7056000
X420 24 395 inv02 $T=3705000 7056000 1 180 $X=3680000 $Y=7056000
X421 24 396 inv02 $T=3696000 10304000 0 0 $X=3696000 $Y=10304000
X422 24 397 inv02 $T=3696000 12624000 0 0 $X=3696000 $Y=12624000
X423 24 398 inv02 $T=3737000 7520000 1 180 $X=3712000 $Y=7520000
X424 24 399 inv02 $T=3728000 6128000 0 0 $X=3728000 $Y=6128000
X425 24 400 inv02 $T=3728000 10304000 0 0 $X=3728000 $Y=10304000
X426 24 401 inv02 $T=3753000 12624000 1 180 $X=3728000 $Y=12624000
X427 24 402 inv02 $T=3744000 7520000 0 0 $X=3744000 $Y=7520000
X428 24 403 inv02 $T=3769000 11928000 1 180 $X=3744000 $Y=11928000
X429 24 404 inv02 $T=3752000 2416000 0 0 $X=3752000 $Y=2416000
X430 24 405 inv02 $T=3816000 10304000 0 0 $X=3816000 $Y=10304000
X431 24 406 inv02 $T=3840000 5432000 0 0 $X=3840000 $Y=5432000
X432 24 407 inv02 $T=4041000 7056000 1 180 $X=4016000 $Y=7056000
X433 24 408 inv02 $T=4041000 11696000 1 180 $X=4016000 $Y=11696000
X434 24 409 inv02 $T=4032000 10072000 0 0 $X=4032000 $Y=10072000
X435 24 410 inv02 $T=4065000 6360000 1 180 $X=4040000 $Y=6360000
X436 24 411 inv02 $T=4040000 11232000 0 0 $X=4040000 $Y=11232000
X437 24 412 inv02 $T=4089000 6128000 1 180 $X=4064000 $Y=6128000
X438 24 413 inv02 $T=4072000 6360000 0 0 $X=4072000 $Y=6360000
X439 24 414 inv02 $T=4096000 6128000 0 0 $X=4096000 $Y=6128000
X440 24 415 inv02 $T=4145000 11928000 1 180 $X=4120000 $Y=11928000
X441 24 416 inv02 $T=4152000 6824000 0 0 $X=4152000 $Y=6824000
X442 24 417 inv02 $T=4200000 12624000 0 0 $X=4200000 $Y=12624000
X443 24 418 inv02 $T=4297000 12624000 1 180 $X=4272000 $Y=12624000
X444 24 419 inv02 $T=4304000 8448000 0 0 $X=4304000 $Y=8448000
X445 24 420 inv02 $T=4304000 9840000 0 0 $X=4304000 $Y=9840000
X446 24 421 inv02 $T=4304000 12624000 0 0 $X=4304000 $Y=12624000
X447 24 422 inv02 $T=4337000 7984000 1 180 $X=4312000 $Y=7984000
X448 24 423 inv02 $T=4345000 9376000 1 180 $X=4320000 $Y=9376000
X449 24 424 inv02 $T=4336000 11000000 0 0 $X=4336000 $Y=11000000
X450 24 425 inv02 $T=4336000 12624000 0 0 $X=4336000 $Y=12624000
X451 24 426 inv02 $T=4344000 4040000 0 0 $X=4344000 $Y=4040000
X452 24 427 inv02 $T=4377000 7288000 1 180 $X=4352000 $Y=7288000
X453 24 428 inv02 $T=4352000 9376000 0 0 $X=4352000 $Y=9376000
X454 24 429 inv02 $T=4360000 12160000 0 0 $X=4360000 $Y=12160000
X455 24 430 inv02 $T=4385000 12392000 1 180 $X=4360000 $Y=12392000
X456 24 431 inv02 $T=4368000 10768000 0 0 $X=4368000 $Y=10768000
X457 24 432 inv02 $T=4393000 12624000 1 180 $X=4368000 $Y=12624000
X458 24 433 inv02 $T=4392000 9840000 0 0 $X=4392000 $Y=9840000
X459 24 434 inv02 $T=4425000 12624000 1 180 $X=4400000 $Y=12624000
X460 24 435 inv02 $T=4408000 4736000 0 0 $X=4408000 $Y=4736000
X461 24 436 inv02 $T=4424000 2416000 0 0 $X=4424000 $Y=2416000
X462 24 437 inv02 $T=4449000 2648000 1 180 $X=4424000 $Y=2648000
X463 24 438 inv02 $T=4449000 5200000 1 180 $X=4424000 $Y=5200000
X464 24 439 inv02 $T=4432000 12624000 0 0 $X=4432000 $Y=12624000
X465 24 440 inv02 $T=4440000 11928000 0 0 $X=4440000 $Y=11928000
X466 24 441 inv02 $T=4448000 12856000 0 0 $X=4448000 $Y=12856000
X467 24 442 inv02 $T=4489000 12624000 1 180 $X=4464000 $Y=12624000
X468 24 443 inv02 $T=4497000 5896000 1 180 $X=4472000 $Y=5896000
X469 24 444 inv02 $T=4497000 9144000 1 180 $X=4472000 $Y=9144000
X470 24 445 inv02 $T=4497000 12392000 1 180 $X=4472000 $Y=12392000
X471 24 446 inv02 $T=4521000 12624000 1 180 $X=4496000 $Y=12624000
X472 24 447 inv02 $T=4529000 6128000 1 180 $X=4504000 $Y=6128000
X473 24 448 inv02 $T=4593000 10536000 1 180 $X=4568000 $Y=10536000
X474 24 449 inv02 $T=4609000 7752000 1 180 $X=4584000 $Y=7752000
X475 24 450 inv02 $T=4584000 12160000 0 0 $X=4584000 $Y=12160000
X476 24 451 inv02 $T=4600000 6128000 0 0 $X=4600000 $Y=6128000
X477 24 452 inv02 $T=4625000 10536000 1 180 $X=4600000 $Y=10536000
X478 24 453 inv02 $T=4641000 7752000 1 180 $X=4616000 $Y=7752000
X479 24 454 inv02 $T=4657000 6128000 1 180 $X=4632000 $Y=6128000
X480 24 455 inv02 $T=4632000 9376000 0 0 $X=4632000 $Y=9376000
X481 24 456 inv02 $T=4681000 7056000 1 180 $X=4656000 $Y=7056000
X482 24 457 inv02 $T=4689000 6128000 1 180 $X=4664000 $Y=6128000
X483 24 458 inv02 $T=4689000 8216000 1 180 $X=4664000 $Y=8216000
X484 24 459 inv02 $T=4688000 11696000 0 0 $X=4688000 $Y=11696000
X485 24 460 inv02 $T=4696000 6128000 0 0 $X=4696000 $Y=6128000
X486 24 461 inv02 $T=4745000 4040000 1 180 $X=4720000 $Y=4040000
X487 24 462 inv02 $T=4745000 10304000 1 180 $X=4720000 $Y=10304000
X488 24 463 inv02 $T=4728000 6128000 0 0 $X=4728000 $Y=6128000
X489 24 464 inv02 $T=4761000 8680000 1 180 $X=4736000 $Y=8680000
X490 24 465 inv02 $T=4736000 8912000 0 0 $X=4736000 $Y=8912000
X491 24 466 inv02 $T=4752000 4040000 0 0 $X=4752000 $Y=4040000
X492 24 467 inv02 $T=4752000 5896000 0 0 $X=4752000 $Y=5896000
X493 24 468 inv02 $T=4777000 13088000 1 180 $X=4752000 $Y=13088000
X494 24 469 inv02 $T=4785000 6128000 1 180 $X=4760000 $Y=6128000
X495 24 470 inv02 $T=4793000 5664000 1 180 $X=4768000 $Y=5664000
X496 24 471 inv02 $T=4776000 8216000 0 0 $X=4776000 $Y=8216000
X497 24 472 inv02 $T=4809000 13088000 1 180 $X=4784000 $Y=13088000
X498 24 473 inv02 $T=4792000 6128000 0 0 $X=4792000 $Y=6128000
X499 24 474 inv02 $T=4800000 4736000 0 0 $X=4800000 $Y=4736000
X500 24 475 inv02 $T=4825000 5664000 1 180 $X=4800000 $Y=5664000
X501 24 476 inv02 $T=4825000 10536000 1 180 $X=4800000 $Y=10536000
X502 24 477 inv02 $T=4816000 13088000 0 0 $X=4816000 $Y=13088000
X503 24 478 inv02 $T=4824000 6128000 0 0 $X=4824000 $Y=6128000
X504 24 479 inv02 $T=4849000 11696000 1 180 $X=4824000 $Y=11696000
X505 24 480 inv02 $T=4857000 5664000 1 180 $X=4832000 $Y=5664000
X506 24 481 inv02 $T=4865000 7984000 1 180 $X=4840000 $Y=7984000
X507 24 482 inv02 $T=4881000 6128000 1 180 $X=4856000 $Y=6128000
X508 24 483 inv02 $T=4889000 5664000 1 180 $X=4864000 $Y=5664000
X509 24 484 inv02 $T=4888000 6128000 0 0 $X=4888000 $Y=6128000
X510 24 485 inv02 $T=4904000 11928000 0 0 $X=4904000 $Y=11928000
X511 24 486 inv02 $T=4945000 6128000 1 180 $X=4920000 $Y=6128000
X512 24 487 inv02 $T=4976000 12160000 0 0 $X=4976000 $Y=12160000
X513 24 488 inv02 $T=5008000 10304000 0 0 $X=5008000 $Y=10304000
X514 24 489 inv02 $T=5032000 9376000 0 0 $X=5032000 $Y=9376000
X515 24 490 inv02 $T=5040000 7752000 0 0 $X=5040000 $Y=7752000
X516 24 491 inv02 $T=5048000 9608000 0 0 $X=5048000 $Y=9608000
X517 24 492 inv02 $T=5089000 1720000 1 180 $X=5064000 $Y=1720000
X518 24 493 inv02 $T=5121000 4272000 1 180 $X=5096000 $Y=4272000
X519 24 494 inv02 $T=5121000 10304000 1 180 $X=5096000 $Y=10304000
X520 24 495 inv02 $T=5120000 8912000 0 0 $X=5120000 $Y=8912000
X521 24 496 inv02 $T=5120000 10536000 0 0 $X=5120000 $Y=10536000
X522 24 497 inv02 $T=5208000 11000000 0 0 $X=5208000 $Y=11000000
X523 24 498 inv02 $T=5216000 12392000 0 0 $X=5216000 $Y=12392000
X524 24 499 inv02 $T=5224000 12160000 0 0 $X=5224000 $Y=12160000
X525 24 500 inv02 $T=5232000 12624000 0 0 $X=5232000 $Y=12624000
X526 24 501 inv02 $T=5265000 9144000 1 180 $X=5240000 $Y=9144000
X527 24 502 inv02 $T=5248000 10072000 0 0 $X=5248000 $Y=10072000
X528 24 503 inv02 $T=5264000 12624000 0 0 $X=5264000 $Y=12624000
X529 24 504 inv02 $T=5305000 11000000 1 180 $X=5280000 $Y=11000000
X530 24 505 inv02 $T=5296000 12624000 0 0 $X=5296000 $Y=12624000
X531 24 506 inv02 $T=5328000 11232000 0 0 $X=5328000 $Y=11232000
X532 24 507 inv02 $T=5352000 560000 0 0 $X=5352000 $Y=560000
X533 24 508 inv02 $T=5360000 9608000 0 0 $X=5360000 $Y=9608000
X534 24 509 inv02 $T=5400000 13088000 0 0 $X=5400000 $Y=13088000
X535 24 510 inv02 $T=5416000 96000 0 0 $X=5416000 $Y=96000
X536 24 511 inv02 $T=5497000 328000 1 180 $X=5472000 $Y=328000
X537 24 512 inv02 $T=5497000 8448000 1 180 $X=5472000 $Y=8448000
X538 24 513 inv02 $T=5472000 10304000 0 0 $X=5472000 $Y=10304000
X539 24 514 inv02 $T=5529000 8448000 1 180 $X=5504000 $Y=8448000
X540 24 515 inv02 $T=5561000 8448000 1 180 $X=5536000 $Y=8448000
X541 24 516 inv02 $T=5593000 8448000 1 180 $X=5568000 $Y=8448000
X542 24 517 inv02 $T=5617000 11696000 1 180 $X=5592000 $Y=11696000
X543 24 518 inv02 $T=5625000 7752000 1 180 $X=5600000 $Y=7752000
X544 24 519 inv02 $T=5625000 8448000 1 180 $X=5600000 $Y=8448000
X545 24 520 inv02 $T=5633000 11232000 1 180 $X=5608000 $Y=11232000
X546 24 521 inv02 $T=5641000 7984000 1 180 $X=5616000 $Y=7984000
X547 24 522 inv02 $T=5624000 7520000 0 0 $X=5624000 $Y=7520000
X548 24 523 inv02 $T=5624000 9840000 0 0 $X=5624000 $Y=9840000
X549 24 524 inv02 $T=5657000 8448000 1 180 $X=5632000 $Y=8448000
X550 24 525 inv02 $T=5640000 3808000 0 0 $X=5640000 $Y=3808000
X551 24 526 inv02 $T=5640000 11232000 0 0 $X=5640000 $Y=11232000
X552 24 527 inv02 $T=5656000 8680000 0 0 $X=5656000 $Y=8680000
X553 24 528 inv02 $T=5681000 9840000 1 180 $X=5656000 $Y=9840000
X554 24 529 inv02 $T=5672000 3808000 0 0 $X=5672000 $Y=3808000
X555 24 530 inv02 $T=5680000 9376000 0 0 $X=5680000 $Y=9376000
X556 24 531 inv02 $T=5729000 8448000 1 180 $X=5704000 $Y=8448000
X557 24 532 inv02 $T=5712000 11000000 0 0 $X=5712000 $Y=11000000
X558 24 533 inv02 $T=5753000 12624000 1 180 $X=5728000 $Y=12624000
X559 24 534 inv02 $T=5736000 8448000 0 0 $X=5736000 $Y=8448000
X560 24 535 inv02 $T=5768000 9144000 0 0 $X=5768000 $Y=9144000
X561 24 536 inv02 $T=5825000 11000000 1 180 $X=5800000 $Y=11000000
X562 24 537 inv02 $T=5808000 8448000 0 0 $X=5808000 $Y=8448000
X563 24 538 inv02 $T=5808000 9840000 0 0 $X=5808000 $Y=9840000
X564 24 539 inv02 $T=5833000 10536000 1 180 $X=5808000 $Y=10536000
X565 24 540 inv02 $T=5840000 3112000 0 0 $X=5840000 $Y=3112000
X566 24 541 inv02 $T=5840000 8448000 0 0 $X=5840000 $Y=8448000
X567 24 542 inv02 $T=5840000 13320000 0 0 $X=5840000 $Y=13320000
X568 24 543 inv02 $T=5848000 11232000 0 0 $X=5848000 $Y=11232000
X569 24 544 inv02 $T=5881000 12624000 1 180 $X=5856000 $Y=12624000
X570 24 545 inv02 $T=5897000 3112000 1 180 $X=5872000 $Y=3112000
X571 24 546 inv02 $T=5872000 8912000 0 0 $X=5872000 $Y=8912000
X572 24 547 inv02 $T=5905000 4736000 1 180 $X=5880000 $Y=4736000
X573 24 548 inv02 $T=5905000 11232000 1 180 $X=5880000 $Y=11232000
X574 24 549 inv02 $T=5888000 12624000 0 0 $X=5888000 $Y=12624000
X575 24 550 inv02 $T=5904000 3112000 0 0 $X=5904000 $Y=3112000
X576 24 551 inv02 $T=5937000 13320000 1 180 $X=5912000 $Y=13320000
X577 24 552 inv02 $T=5945000 2648000 1 180 $X=5920000 $Y=2648000
X578 24 553 inv02 $T=5920000 12624000 0 0 $X=5920000 $Y=12624000
X579 24 554 inv02 $T=5945000 12856000 1 180 $X=5920000 $Y=12856000
X580 24 555 inv02 $T=5961000 7984000 1 180 $X=5936000 $Y=7984000
X581 24 556 inv02 $T=5961000 11464000 1 180 $X=5936000 $Y=11464000
X582 24 557 inv02 $T=5944000 2880000 0 0 $X=5944000 $Y=2880000
X583 24 558 inv02 $T=5944000 13320000 0 0 $X=5944000 $Y=13320000
X584 24 559 inv02 $T=5977000 2648000 1 180 $X=5952000 $Y=2648000
X585 24 560 inv02 $T=5977000 4272000 1 180 $X=5952000 $Y=4272000
X586 24 561 inv02 $T=5977000 12624000 1 180 $X=5952000 $Y=12624000
X587 24 562 inv02 $T=5952000 12856000 0 0 $X=5952000 $Y=12856000
X588 24 563 inv02 $T=5985000 8912000 1 180 $X=5960000 $Y=8912000
X589 24 564 inv02 $T=5960000 11928000 0 0 $X=5960000 $Y=11928000
X590 24 565 inv02 $T=5968000 8216000 0 0 $X=5968000 $Y=8216000
X591 24 566 inv02 $T=5993000 11232000 1 180 $X=5968000 $Y=11232000
X592 24 567 inv02 $T=5993000 11464000 1 180 $X=5968000 $Y=11464000
X593 24 568 inv02 $T=5992000 7752000 0 0 $X=5992000 $Y=7752000
X594 24 569 inv02 $T=6025000 5200000 1 180 $X=6000000 $Y=5200000
X595 24 570 inv02 $T=6024000 7752000 0 0 $X=6024000 $Y=7752000
X596 24 571 inv02 $T=6032000 1024000 0 0 $X=6032000 $Y=1024000
X597 24 572 inv02 $T=6048000 12856000 0 0 $X=6048000 $Y=12856000
X598 24 573 inv02 $T=6113000 7984000 1 180 $X=6088000 $Y=7984000
X599 24 574 inv02 $T=6113000 9376000 1 180 $X=6088000 $Y=9376000
X600 24 575 inv02 $T=6113000 10536000 1 180 $X=6088000 $Y=10536000
X601 24 576 inv02 $T=6121000 12624000 1 180 $X=6096000 $Y=12624000
X602 24 577 inv02 $T=6137000 7752000 1 180 $X=6112000 $Y=7752000
X603 24 578 inv02 $T=6145000 6824000 1 180 $X=6120000 $Y=6824000
X604 24 579 inv02 $T=6120000 9376000 0 0 $X=6120000 $Y=9376000
X605 24 580 inv02 $T=6169000 7752000 1 180 $X=6144000 $Y=7752000
X606 24 581 inv02 $T=6184000 328000 0 0 $X=6184000 $Y=328000
X607 24 582 inv02 $T=6216000 328000 0 0 $X=6216000 $Y=328000
X608 24 583 inv02 $T=6257000 5432000 1 180 $X=6232000 $Y=5432000
X609 24 584 inv02 $T=6257000 8448000 1 180 $X=6232000 $Y=8448000
X610 24 585 inv02 $T=6248000 9840000 0 0 $X=6248000 $Y=9840000
X611 24 586 inv02 $T=6289000 2648000 1 180 $X=6264000 $Y=2648000
X612 24 587 inv02 $T=6304000 8448000 0 0 $X=6304000 $Y=8448000
X613 24 588 inv02 $T=6337000 2880000 1 180 $X=6312000 $Y=2880000
X614 24 589 inv02 $T=6345000 6360000 1 180 $X=6320000 $Y=6360000
X615 24 590 inv02 $T=6320000 9840000 0 0 $X=6320000 $Y=9840000
X616 24 591 inv02 $T=6320000 13320000 0 0 $X=6320000 $Y=13320000
X617 24 592 inv02 $T=6353000 1488000 1 180 $X=6328000 $Y=1488000
X618 24 593 inv02 $T=6336000 7984000 0 0 $X=6336000 $Y=7984000
X619 24 594 inv02 $T=6369000 1024000 1 180 $X=6344000 $Y=1024000
X620 24 595 inv02 $T=6377000 6360000 1 180 $X=6352000 $Y=6360000
X621 24 596 inv02 $T=6377000 9840000 1 180 $X=6352000 $Y=9840000
X622 24 597 inv02 $T=6368000 12160000 0 0 $X=6368000 $Y=12160000
X623 24 598 inv02 $T=6401000 3344000 1 180 $X=6376000 $Y=3344000
X624 24 599 inv02 $T=6401000 9144000 1 180 $X=6376000 $Y=9144000
X625 24 600 inv02 $T=6376000 10072000 0 0 $X=6376000 $Y=10072000
X626 24 601 inv02 $T=6409000 560000 1 180 $X=6384000 $Y=560000
X627 24 602 inv02 $T=6384000 792000 0 0 $X=6384000 $Y=792000
X628 24 603 inv02 $T=6384000 2416000 0 0 $X=6384000 $Y=2416000
X629 24 604 inv02 $T=6400000 8912000 0 0 $X=6400000 $Y=8912000
X630 24 605 inv02 $T=6400000 12160000 0 0 $X=6400000 $Y=12160000
X631 24 606 inv02 $T=6433000 3344000 1 180 $X=6408000 $Y=3344000
X632 24 607 inv02 $T=6408000 12392000 0 0 $X=6408000 $Y=12392000
X633 24 608 inv02 $T=6433000 12624000 1 180 $X=6408000 $Y=12624000
X634 24 609 inv02 $T=6449000 7752000 1 180 $X=6424000 $Y=7752000
X635 24 610 inv02 $T=6432000 8912000 0 0 $X=6432000 $Y=8912000
X636 24 611 inv02 $T=6432000 12160000 0 0 $X=6432000 $Y=12160000
X637 24 612 inv02 $T=6440000 9376000 0 0 $X=6440000 $Y=9376000
X638 24 613 inv02 $T=6465000 12392000 1 180 $X=6440000 $Y=12392000
X639 24 614 inv02 $T=6489000 6824000 1 180 $X=6464000 $Y=6824000
X640 24 615 inv02 $T=6489000 8912000 1 180 $X=6464000 $Y=8912000
X641 24 616 inv02 $T=6464000 12160000 0 0 $X=6464000 $Y=12160000
X642 24 617 inv02 $T=6497000 9376000 1 180 $X=6472000 $Y=9376000
X643 24 618 inv02 $T=6497000 12392000 1 180 $X=6472000 $Y=12392000
X644 24 619 inv02 $T=6488000 8680000 0 0 $X=6488000 $Y=8680000
X645 24 620 inv02 $T=6521000 6824000 1 180 $X=6496000 $Y=6824000
X646 24 621 inv02 $T=6496000 8216000 0 0 $X=6496000 $Y=8216000
X647 24 622 inv02 $T=6496000 8912000 0 0 $X=6496000 $Y=8912000
X648 24 623 inv02 $T=6521000 12160000 1 180 $X=6496000 $Y=12160000
X649 24 624 inv02 $T=6529000 12392000 1 180 $X=6504000 $Y=12392000
X650 24 625 inv02 $T=6545000 8680000 1 180 $X=6520000 $Y=8680000
X651 24 626 inv02 $T=6552000 8680000 0 0 $X=6552000 $Y=8680000
X652 24 627 inv02 $T=6609000 8680000 1 180 $X=6584000 $Y=8680000
X653 24 628 inv02 $T=6616000 5896000 0 0 $X=6616000 $Y=5896000
X654 24 629 inv02 $T=6616000 8680000 0 0 $X=6616000 $Y=8680000
X655 24 630 inv02 $T=6649000 96000 1 180 $X=6624000 $Y=96000
X656 24 631 inv02 $T=6648000 8680000 0 0 $X=6648000 $Y=8680000
X657 24 632 inv02 $T=6648000 11928000 0 0 $X=6648000 $Y=11928000
X658 24 633 inv02 $T=6705000 11928000 1 180 $X=6680000 $Y=11928000
X659 24 634 inv02 $T=6721000 6360000 1 180 $X=6696000 $Y=6360000
X660 24 635 inv02 $T=6696000 10072000 0 0 $X=6696000 $Y=10072000
X661 24 636 inv02 $T=6712000 11928000 0 0 $X=6712000 $Y=11928000
X662 24 637 inv02 $T=6736000 1720000 0 0 $X=6736000 $Y=1720000
X663 24 638 inv02 $T=6744000 11928000 0 0 $X=6744000 $Y=11928000
X664 24 639 inv02 $T=6849000 12160000 1 180 $X=6824000 $Y=12160000
X665 24 640 inv02 $T=6848000 1024000 0 0 $X=6848000 $Y=1024000
X666 24 641 inv02 $T=6848000 11232000 0 0 $X=6848000 $Y=11232000
X667 24 642 inv02 $T=6856000 328000 0 0 $X=6856000 $Y=328000
X668 24 643 inv02 $T=6856000 12160000 0 0 $X=6856000 $Y=12160000
X669 24 644 inv02 $T=6913000 4272000 1 180 $X=6888000 $Y=4272000
X670 24 645 inv02 $T=6921000 11000000 1 180 $X=6896000 $Y=11000000
X671 24 646 inv02 $T=6904000 11464000 0 0 $X=6904000 $Y=11464000
X672 24 647 inv02 $T=6937000 5432000 1 180 $X=6912000 $Y=5432000
X673 24 648 inv02 $T=6945000 4272000 1 180 $X=6920000 $Y=4272000
X674 24 649 inv02 $T=6953000 11000000 1 180 $X=6928000 $Y=11000000
X675 24 650 inv02 $T=6961000 11464000 1 180 $X=6936000 $Y=11464000
X676 24 651 inv02 $T=6969000 13320000 1 180 $X=6944000 $Y=13320000
X677 24 652 inv02 $T=6977000 4272000 1 180 $X=6952000 $Y=4272000
X678 24 653 inv02 $T=6977000 12160000 1 180 $X=6952000 $Y=12160000
X679 24 654 inv02 $T=6993000 11464000 1 180 $X=6968000 $Y=11464000
X680 24 655 inv02 $T=7001000 6360000 1 180 $X=6976000 $Y=6360000
X681 24 656 inv02 $T=7009000 12160000 1 180 $X=6984000 $Y=12160000
X682 24 657 inv02 $T=7041000 3112000 1 180 $X=7016000 $Y=3112000
X683 24 658 inv02 $T=7024000 11928000 0 0 $X=7024000 $Y=11928000
X684 24 659 inv02 $T=7048000 3112000 0 0 $X=7048000 $Y=3112000
X685 24 660 inv02 $T=7080000 3112000 0 0 $X=7080000 $Y=3112000
X686 24 661 inv02 $T=7185000 4504000 1 180 $X=7160000 $Y=4504000
X687 24 662 inv02 $T=7201000 3112000 1 180 $X=7176000 $Y=3112000
X688 24 663 inv02 $T=7209000 12160000 1 180 $X=7184000 $Y=12160000
X689 24 664 inv02 $T=7192000 4504000 0 0 $X=7192000 $Y=4504000
X690 24 665 inv02 $T=7233000 96000 1 180 $X=7208000 $Y=96000
X691 24 666 inv02 $T=7265000 11232000 1 180 $X=7240000 $Y=11232000
X692 24 667 inv02 $T=7256000 13320000 0 0 $X=7256000 $Y=13320000
X693 24 668 inv02 $T=7297000 11232000 1 180 $X=7272000 $Y=11232000
X694 24 669 inv02 $T=7313000 10768000 1 180 $X=7288000 $Y=10768000
X695 24 670 inv02 $T=7313000 13320000 1 180 $X=7288000 $Y=13320000
X696 24 671 inv02 $T=7321000 11000000 1 180 $X=7296000 $Y=11000000
X697 24 672 inv02 $T=7304000 12624000 0 0 $X=7304000 $Y=12624000
X698 24 673 inv02 $T=7320000 10768000 0 0 $X=7320000 $Y=10768000
X699 24 674 inv02 $T=7328000 2416000 0 0 $X=7328000 $Y=2416000
X700 24 675 inv02 $T=7336000 12624000 0 0 $X=7336000 $Y=12624000
X701 24 676 inv02 $T=7344000 11232000 0 0 $X=7344000 $Y=11232000
X702 24 677 inv02 $T=7360000 2416000 0 0 $X=7360000 $Y=2416000
X703 24 678 inv02 $T=7368000 12624000 0 0 $X=7368000 $Y=12624000
X704 24 679 inv02 $T=7401000 4040000 1 180 $X=7376000 $Y=4040000
X705 24 680 inv02 $T=7376000 11232000 0 0 $X=7376000 $Y=11232000
X706 24 681 inv02 $T=7392000 1024000 0 0 $X=7392000 $Y=1024000
X707 24 682 inv02 $T=7392000 5664000 0 0 $X=7392000 $Y=5664000
X708 24 683 inv02 $T=7392000 7056000 0 0 $X=7392000 $Y=7056000
X709 24 684 inv02 $T=7441000 11928000 1 180 $X=7416000 $Y=11928000
X710 24 685 inv02 $T=7424000 5664000 0 0 $X=7424000 $Y=5664000
X711 24 686 inv02 $T=7432000 328000 0 0 $X=7432000 $Y=328000
X712 24 687 inv02 $T=7448000 3344000 0 0 $X=7448000 $Y=3344000
X713 24 688 inv02 $T=7464000 328000 0 0 $X=7464000 $Y=328000
X714 24 689 inv02 $T=7489000 4040000 1 180 $X=7464000 $Y=4040000
X715 24 690 inv02 $T=7521000 9608000 1 180 $X=7496000 $Y=9608000
X716 24 691 inv02 $T=7529000 9376000 1 180 $X=7504000 $Y=9376000
X717 24 692 inv02 $T=7537000 12160000 1 180 $X=7512000 $Y=12160000
X718 24 693 inv02 $T=7536000 9376000 0 0 $X=7536000 $Y=9376000
X719 24 694 inv02 $T=7585000 328000 1 180 $X=7560000 $Y=328000
X720 24 695 inv02 $T=7593000 9376000 1 180 $X=7568000 $Y=9376000
X721 24 696 inv02 $T=7641000 8680000 1 180 $X=7616000 $Y=8680000
X722 24 697 inv02 $T=7632000 3808000 0 0 $X=7632000 $Y=3808000
X723 24 698 inv02 $T=7648000 8680000 0 0 $X=7648000 $Y=8680000
X724 24 699 inv02 $T=7672000 7056000 0 0 $X=7672000 $Y=7056000
X725 24 700 inv02 $T=7721000 4968000 1 180 $X=7696000 $Y=4968000
X726 24 701 inv02 $T=7737000 12392000 1 180 $X=7712000 $Y=12392000
X727 24 702 inv02 $T=7744000 12392000 0 0 $X=7744000 $Y=12392000
X728 24 703 inv02 $T=7752000 11928000 0 0 $X=7752000 $Y=11928000
X729 24 704 inv02 $T=7776000 12392000 0 0 $X=7776000 $Y=12392000
X730 24 705 inv02 $T=7817000 3112000 1 180 $X=7792000 $Y=3112000
X731 24 706 inv02 $T=7800000 12856000 0 0 $X=7800000 $Y=12856000
X732 24 707 inv02 $T=7833000 560000 1 180 $X=7808000 $Y=560000
X733 24 708 inv02 $T=7833000 9608000 1 180 $X=7808000 $Y=9608000
X734 24 709 inv02 $T=7833000 12392000 1 180 $X=7808000 $Y=12392000
X735 24 710 inv02 $T=7824000 3112000 0 0 $X=7824000 $Y=3112000
X736 24 711 inv02 $T=7840000 560000 0 0 $X=7840000 $Y=560000
X737 24 712 inv02 $T=7865000 9608000 1 180 $X=7840000 $Y=9608000
X738 24 713 inv02 $T=7840000 12392000 0 0 $X=7840000 $Y=12392000
X739 24 714 inv02 $T=7848000 10072000 0 0 $X=7848000 $Y=10072000
X740 24 715 inv02 $T=7848000 12160000 0 0 $X=7848000 $Y=12160000
X741 24 716 inv02 $T=7897000 9608000 1 180 $X=7872000 $Y=9608000
X742 24 717 inv02 $T=7872000 12392000 0 0 $X=7872000 $Y=12392000
X743 24 718 inv02 $T=7905000 4272000 1 180 $X=7880000 $Y=4272000
X744 24 719 inv02 $T=7880000 10072000 0 0 $X=7880000 $Y=10072000
X745 24 720 inv02 $T=7880000 12160000 0 0 $X=7880000 $Y=12160000
X746 24 721 inv02 $T=7904000 9144000 0 0 $X=7904000 $Y=9144000
X747 24 722 inv02 $T=7929000 9608000 1 180 $X=7904000 $Y=9608000
X748 24 723 inv02 $T=7904000 12392000 0 0 $X=7904000 $Y=12392000
X749 24 724 inv02 $T=7937000 10072000 1 180 $X=7912000 $Y=10072000
X750 24 725 inv02 $T=7936000 1488000 0 0 $X=7936000 $Y=1488000
X751 24 726 inv02 $T=7936000 9144000 0 0 $X=7936000 $Y=9144000
X752 24 727 inv02 $T=7961000 12392000 1 180 $X=7936000 $Y=12392000
X753 24 728 inv02 $T=7969000 10072000 1 180 $X=7944000 $Y=10072000
X754 24 729 inv02 $T=7960000 8680000 0 0 $X=7960000 $Y=8680000
X755 24 730 inv02 $T=7968000 1488000 0 0 $X=7968000 $Y=1488000
X756 24 731 inv02 $T=7993000 2880000 1 180 $X=7968000 $Y=2880000
X757 24 732 inv02 $T=7993000 12392000 1 180 $X=7968000 $Y=12392000
X758 24 733 inv02 $T=8001000 10072000 1 180 $X=7976000 $Y=10072000
X759 24 734 inv02 $T=7984000 8912000 0 0 $X=7984000 $Y=8912000
X760 24 735 inv02 $T=7992000 8680000 0 0 $X=7992000 $Y=8680000
X761 24 736 inv02 $T=8000000 1488000 0 0 $X=8000000 $Y=1488000
X762 24 737 inv02 $T=8000000 2880000 0 0 $X=8000000 $Y=2880000
X763 24 738 inv02 $T=8008000 10072000 0 0 $X=8008000 $Y=10072000
X764 24 739 inv02 $T=8041000 8912000 1 180 $X=8016000 $Y=8912000
X765 24 740 inv02 $T=8024000 4040000 0 0 $X=8024000 $Y=4040000
X766 24 741 inv02 $T=8024000 5896000 0 0 $X=8024000 $Y=5896000
X767 24 742 inv02 $T=8032000 1488000 0 0 $X=8032000 $Y=1488000
X768 24 743 inv02 $T=8057000 7984000 1 180 $X=8032000 $Y=7984000
X769 24 744 inv02 $T=8057000 8216000 1 180 $X=8032000 $Y=8216000
X770 24 745 inv02 $T=8040000 10072000 0 0 $X=8040000 $Y=10072000
X771 24 746 inv02 $T=8048000 6128000 0 0 $X=8048000 $Y=6128000
X772 24 747 inv02 $T=8073000 8912000 1 180 $X=8048000 $Y=8912000
X773 24 748 inv02 $T=8056000 4040000 0 0 $X=8056000 $Y=4040000
X774 24 749 inv02 $T=8056000 5896000 0 0 $X=8056000 $Y=5896000
X775 24 750 inv02 $T=8089000 8216000 1 180 $X=8064000 $Y=8216000
X776 24 751 inv02 $T=8072000 792000 0 0 $X=8072000 $Y=792000
X777 24 752 inv02 $T=8088000 4040000 0 0 $X=8088000 $Y=4040000
X778 24 753 inv02 $T=8096000 8216000 0 0 $X=8096000 $Y=8216000
X779 24 754 inv02 $T=8120000 4040000 0 0 $X=8120000 $Y=4040000
X780 24 755 inv02 $T=8128000 8216000 0 0 $X=8128000 $Y=8216000
X781 24 756 inv02 $T=8136000 1024000 0 0 $X=8136000 $Y=1024000
X782 24 757 inv02 $T=8177000 4040000 1 180 $X=8152000 $Y=4040000
X783 24 758 inv02 $T=8200000 5200000 0 0 $X=8200000 $Y=5200000
X784 24 759 inv02 $T=8225000 13088000 1 180 $X=8200000 $Y=13088000
X785 24 760 inv02 $T=8216000 792000 0 0 $X=8216000 $Y=792000
X786 24 761 inv02 $T=8216000 3808000 0 0 $X=8216000 $Y=3808000
X787 24 762 inv02 $T=8241000 9144000 1 180 $X=8216000 $Y=9144000
X788 24 763 inv02 $T=8257000 560000 1 180 $X=8232000 $Y=560000
X789 24 764 inv02 $T=8232000 5200000 0 0 $X=8232000 $Y=5200000
X790 24 765 inv02 $T=8248000 9144000 0 0 $X=8248000 $Y=9144000
X791 24 766 inv02 $T=8297000 8680000 1 180 $X=8272000 $Y=8680000
X792 24 767 inv02 $T=8352000 8680000 0 0 $X=8352000 $Y=8680000
X793 24 768 inv02 $T=8368000 7752000 0 0 $X=8368000 $Y=7752000
X794 24 769 inv02 $T=8384000 4968000 0 0 $X=8384000 $Y=4968000
X795 24 770 inv02 $T=8392000 10768000 0 0 $X=8392000 $Y=10768000
X796 24 771 inv02 $T=8425000 7056000 1 180 $X=8400000 $Y=7056000
X797 24 772 inv02 $T=8425000 7752000 1 180 $X=8400000 $Y=7752000
X798 24 773 inv02 $T=8424000 10536000 0 0 $X=8424000 $Y=10536000
X799 24 774 inv02 $T=8432000 5432000 0 0 $X=8432000 $Y=5432000
X800 24 775 inv02 $T=8432000 7056000 0 0 $X=8432000 $Y=7056000
X801 24 776 inv02 $T=8432000 7752000 0 0 $X=8432000 $Y=7752000
X802 24 777 inv02 $T=8473000 1952000 1 180 $X=8448000 $Y=1952000
X803 24 778 inv02 $T=8456000 10536000 0 0 $X=8456000 $Y=10536000
X804 24 779 inv02 $T=8464000 792000 0 0 $X=8464000 $Y=792000
X805 24 780 inv02 $T=8464000 3112000 0 0 $X=8464000 $Y=3112000
X806 24 781 inv02 $T=8464000 4272000 0 0 $X=8464000 $Y=4272000
X807 24 782 inv02 $T=8464000 5432000 0 0 $X=8464000 $Y=5432000
X808 24 783 inv02 $T=8489000 7056000 1 180 $X=8464000 $Y=7056000
X809 24 784 inv02 $T=8480000 6824000 0 0 $X=8480000 $Y=6824000
X810 24 785 inv02 $T=8488000 12160000 0 0 $X=8488000 $Y=12160000
X811 24 786 inv02 $T=8496000 5432000 0 0 $X=8496000 $Y=5432000
X812 24 787 inv02 $T=8496000 7056000 0 0 $X=8496000 $Y=7056000
X813 24 788 inv02 $T=8504000 328000 0 0 $X=8504000 $Y=328000
X814 24 789 inv02 $T=8528000 5432000 0 0 $X=8528000 $Y=5432000
X815 24 790 inv02 $T=8576000 7288000 0 0 $X=8576000 $Y=7288000
X816 24 791 inv02 $T=8576000 9840000 0 0 $X=8576000 $Y=9840000
X817 24 792 inv02 $T=8576000 11928000 0 0 $X=8576000 $Y=11928000
X818 24 793 inv02 $T=8592000 328000 0 0 $X=8592000 $Y=328000
X819 24 794 inv02 $T=8641000 560000 1 180 $X=8616000 $Y=560000
X820 24 795 inv02 $T=8641000 7984000 1 180 $X=8616000 $Y=7984000
X821 24 796 inv02 $T=8649000 328000 1 180 $X=8624000 $Y=328000
X822 24 797 inv02 $T=8673000 560000 1 180 $X=8648000 $Y=560000
X823 24 798 inv02 $T=8648000 2648000 0 0 $X=8648000 $Y=2648000
X824 24 799 inv02 $T=8656000 328000 0 0 $X=8656000 $Y=328000
X825 24 800 inv02 $T=8664000 9840000 0 0 $X=8664000 $Y=9840000
X826 24 801 inv02 $T=8664000 11000000 0 0 $X=8664000 $Y=11000000
X827 24 802 inv02 $T=8689000 13320000 1 180 $X=8664000 $Y=13320000
X828 24 803 inv02 $T=8680000 560000 0 0 $X=8680000 $Y=560000
X829 24 804 inv02 $T=8688000 8912000 0 0 $X=8688000 $Y=8912000
X830 24 805 inv02 $T=8737000 560000 1 180 $X=8712000 $Y=560000
X831 24 806 inv02 $T=8712000 8216000 0 0 $X=8712000 $Y=8216000
X832 24 807 inv02 $T=8745000 8912000 1 180 $X=8720000 $Y=8912000
X833 24 808 inv02 $T=8753000 1952000 1 180 $X=8728000 $Y=1952000
X834 24 809 inv02 $T=8744000 8680000 0 0 $X=8744000 $Y=8680000
X835 24 810 inv02 $T=8752000 328000 0 0 $X=8752000 $Y=328000
X836 24 811 inv02 $T=8752000 8912000 0 0 $X=8752000 $Y=8912000
X837 24 812 inv02 $T=8768000 12160000 0 0 $X=8768000 $Y=12160000
X838 24 813 inv02 $T=8776000 8216000 0 0 $X=8776000 $Y=8216000
X839 24 814 inv02 $T=8776000 8680000 0 0 $X=8776000 $Y=8680000
X840 24 815 inv02 $T=8809000 8912000 1 180 $X=8784000 $Y=8912000
X841 24 816 inv02 $T=8800000 12160000 0 0 $X=8800000 $Y=12160000
X842 24 817 inv02 $T=8857000 7056000 1 180 $X=8832000 $Y=7056000
X843 24 818 inv02 $T=8920000 7288000 0 0 $X=8920000 $Y=7288000
X844 24 819 inv02 $T=8920000 13320000 0 0 $X=8920000 $Y=13320000
X845 24 820 inv02 $T=8977000 7288000 1 180 $X=8952000 $Y=7288000
X846 24 821 inv02 $T=9009000 560000 1 180 $X=8984000 $Y=560000
X847 24 822 inv02 $T=9009000 7288000 1 180 $X=8984000 $Y=7288000
X848 24 823 inv02 $T=8992000 10072000 0 0 $X=8992000 $Y=10072000
X849 24 824 inv02 $T=9025000 11232000 1 180 $X=9000000 $Y=11232000
X850 24 825 inv02 $T=9008000 6824000 0 0 $X=9008000 $Y=6824000
X851 24 826 inv02 $T=9024000 9144000 0 0 $X=9024000 $Y=9144000
X852 24 827 inv02 $T=9049000 10072000 1 180 $X=9024000 $Y=10072000
X853 24 828 inv02 $T=9024000 12624000 0 0 $X=9024000 $Y=12624000
X854 24 829 inv02 $T=9065000 6824000 1 180 $X=9040000 $Y=6824000
X855 24 830 inv02 $T=9081000 8680000 1 180 $X=9056000 $Y=8680000
X856 24 831 inv02 $T=9072000 1952000 0 0 $X=9072000 $Y=1952000
X857 24 832 inv02 $T=9113000 7752000 1 180 $X=9088000 $Y=7752000
X858 24 833 inv02 $T=9096000 10304000 0 0 $X=9096000 $Y=10304000
X859 24 834 inv02 $T=9176000 9840000 0 0 $X=9176000 $Y=9840000
X860 24 835 inv02 $T=9272000 11464000 0 0 $X=9272000 $Y=11464000
X861 24 836 inv02 $T=9320000 6824000 0 0 $X=9320000 $Y=6824000
X862 24 837 inv02 $T=9328000 1256000 0 0 $X=9328000 $Y=1256000
X863 24 838 inv02 $T=9336000 9144000 0 0 $X=9336000 $Y=9144000
X864 24 839 inv02 $T=9416000 11464000 0 0 $X=9416000 $Y=11464000
X865 24 840 inv02 $T=9448000 11464000 0 0 $X=9448000 $Y=11464000
X866 24 841 inv02 $T=9489000 2184000 1 180 $X=9464000 $Y=2184000
X867 24 842 inv02 $T=9489000 9376000 1 180 $X=9464000 $Y=9376000
X868 24 843 inv02 $T=9480000 11464000 0 0 $X=9480000 $Y=11464000
X869 24 844 inv02 $T=9496000 13088000 0 0 $X=9496000 $Y=13088000
X870 24 845 inv02 $T=9537000 11464000 1 180 $X=9512000 $Y=11464000
X871 24 846 inv02 $T=9528000 12160000 0 0 $X=9528000 $Y=12160000
X872 24 847 inv02 $T=9536000 7056000 0 0 $X=9536000 $Y=7056000
X873 24 848 inv02 $T=9560000 12160000 0 0 $X=9560000 $Y=12160000
X874 24 849 inv02 $T=9560000 12392000 0 0 $X=9560000 $Y=12392000
X875 24 850 inv02 $T=9568000 6824000 0 0 $X=9568000 $Y=6824000
X876 24 851 inv02 $T=9617000 3576000 1 180 $X=9592000 $Y=3576000
X877 24 852 inv02 $T=9592000 12160000 0 0 $X=9592000 $Y=12160000
X878 24 853 inv02 $T=9625000 1720000 1 180 $X=9600000 $Y=1720000
X879 24 854 inv02 $T=9625000 6824000 1 180 $X=9600000 $Y=6824000
X880 24 855 inv02 $T=9641000 4504000 1 180 $X=9616000 $Y=4504000
X881 24 856 inv02 $T=9632000 5664000 0 0 $X=9632000 $Y=5664000
X882 24 857 inv02 $T=9632000 6824000 0 0 $X=9632000 $Y=6824000
X883 24 858 inv02 $T=9664000 6824000 0 0 $X=9664000 $Y=6824000
X884 24 859 inv02 $T=9697000 7288000 1 180 $X=9672000 $Y=7288000
X885 24 860 inv02 $T=9721000 6824000 1 180 $X=9696000 $Y=6824000
X886 24 861 inv02 $T=9696000 13552000 0 0 $X=9696000 $Y=13552000
X887 24 862 inv02 $T=9753000 6824000 1 180 $X=9728000 $Y=6824000
X888 24 863 inv02 $T=9760000 6824000 0 0 $X=9760000 $Y=6824000
X889 24 864 inv02 $T=9801000 2184000 1 180 $X=9776000 $Y=2184000
X890 24 865 inv02 $T=9784000 2880000 0 0 $X=9784000 $Y=2880000
X891 24 866 inv02 $T=9792000 6824000 0 0 $X=9792000 $Y=6824000
X892 24 867 inv02 $T=9808000 10768000 0 0 $X=9808000 $Y=10768000
X893 24 868 inv02 $T=9824000 6824000 0 0 $X=9824000 $Y=6824000
X894 24 869 inv02 $T=9840000 4272000 0 0 $X=9840000 $Y=4272000
X895 24 870 inv02 $T=9865000 5200000 1 180 $X=9840000 $Y=5200000
X896 24 871 inv02 $T=9856000 6824000 0 0 $X=9856000 $Y=6824000
X897 24 872 inv02 $T=9905000 12856000 1 180 $X=9880000 $Y=12856000
X898 24 873 inv02 $T=9913000 11464000 1 180 $X=9888000 $Y=11464000
X899 24 874 inv02 $T=9912000 6128000 0 0 $X=9912000 $Y=6128000
X900 24 875 inv02 $T=9937000 12160000 1 180 $X=9912000 $Y=12160000
X901 24 876 inv02 $T=9920000 11464000 0 0 $X=9920000 $Y=11464000
X902 24 877 inv02 $T=9969000 3112000 1 180 $X=9944000 $Y=3112000
X903 24 878 inv02 $T=9944000 12160000 0 0 $X=9944000 $Y=12160000
X904 24 879 inv02 $T=9952000 11696000 0 0 $X=9952000 $Y=11696000
X905 24 880 inv02 $T=9977000 12624000 1 180 $X=9952000 $Y=12624000
X906 24 881 inv02 $T=9993000 12856000 1 180 $X=9968000 $Y=12856000
X907 24 882 inv02 $T=9968000 13088000 0 0 $X=9968000 $Y=13088000
X908 24 883 inv02 $T=9984000 10304000 0 0 $X=9984000 $Y=10304000
X909 24 884 inv02 $T=10080000 12624000 0 0 $X=10080000 $Y=12624000
X910 24 885 inv02 $T=10120000 5200000 0 0 $X=10120000 $Y=5200000
X911 24 886 inv02 $T=10120000 9144000 0 0 $X=10120000 $Y=9144000
X912 24 887 inv02 $T=10177000 2416000 1 180 $X=10152000 $Y=2416000
X913 24 888 inv02 $T=10233000 12856000 1 180 $X=10208000 $Y=12856000
X914 24 889 inv02 $T=10208000 13088000 0 0 $X=10208000 $Y=13088000
X915 24 890 inv02 $T=10232000 5432000 0 0 $X=10232000 $Y=5432000
X916 24 891 inv02 $T=10232000 7752000 0 0 $X=10232000 $Y=7752000
X917 24 892 inv02 $T=10248000 1256000 0 0 $X=10248000 $Y=1256000
X918 24 893 inv02 $T=10296000 12856000 0 0 $X=10296000 $Y=12856000
X919 24 894 inv02 $T=10329000 11928000 1 180 $X=10304000 $Y=11928000
X920 24 895 inv02 $T=10345000 13320000 1 180 $X=10320000 $Y=13320000
X921 24 896 inv02 $T=10336000 792000 0 0 $X=10336000 $Y=792000
X922 24 897 inv02 $T=10360000 11000000 0 0 $X=10360000 $Y=11000000
X923 24 898 inv02 $T=10368000 792000 0 0 $X=10368000 $Y=792000
X924 24 899 inv02 $T=10376000 13088000 0 0 $X=10376000 $Y=13088000
X925 24 900 inv02 $T=10417000 1024000 1 180 $X=10392000 $Y=1024000
X926 24 901 inv02 $T=10400000 2880000 0 0 $X=10400000 $Y=2880000
X927 24 902 inv02 $T=10433000 13088000 1 180 $X=10408000 $Y=13088000
X928 24 903 inv02 $T=10432000 2184000 0 0 $X=10432000 $Y=2184000
X929 24 904 inv02 $T=10432000 10072000 0 0 $X=10432000 $Y=10072000
X930 24 905 inv02 $T=10489000 10072000 1 180 $X=10464000 $Y=10072000
X931 24 906 inv02 $T=10505000 792000 1 180 $X=10480000 $Y=792000
X932 24 907 inv02 $T=10616000 4272000 0 0 $X=10616000 $Y=4272000
X933 24 908 inv02 $T=10648000 4040000 0 0 $X=10648000 $Y=4040000
X934 24 909 inv02 $T=10680000 7984000 0 0 $X=10680000 $Y=7984000
X935 24 910 inv02 $T=10720000 1952000 0 0 $X=10720000 $Y=1952000
X936 24 911 inv02 $T=10785000 7984000 1 180 $X=10760000 $Y=7984000
X937 24 912 inv02 $T=10801000 10072000 1 180 $X=10776000 $Y=10072000
X938 24 913 inv02 $T=10800000 3112000 0 0 $X=10800000 $Y=3112000
X939 24 914 inv02 $T=10833000 10072000 1 180 $X=10808000 $Y=10072000
X940 24 915 inv02 $T=10832000 1024000 0 0 $X=10832000 $Y=1024000
X941 24 916 inv02 $T=10905000 328000 1 180 $X=10880000 $Y=328000
X942 24 917 inv02 $T=10896000 13320000 0 0 $X=10896000 $Y=13320000
X943 24 918 inv02 $T=10953000 11696000 1 180 $X=10928000 $Y=11696000
X944 24 919 inv02 $T=10960000 11696000 0 0 $X=10960000 $Y=11696000
X945 24 920 inv02 $T=10960000 12160000 0 0 $X=10960000 $Y=12160000
X946 24 921 inv02 $T=11049000 792000 1 180 $X=11024000 $Y=792000
X947 24 922 inv02 $T=11048000 13320000 0 0 $X=11048000 $Y=13320000
X948 24 923 inv02 $T=11081000 792000 1 180 $X=11056000 $Y=792000
X949 24 924 inv02 $T=11113000 792000 1 180 $X=11088000 $Y=792000
X950 24 925 inv02 $T=11113000 1488000 1 180 $X=11088000 $Y=1488000
X951 24 926 inv02 $T=11113000 13088000 1 180 $X=11088000 $Y=13088000
X952 24 927 inv02 $T=11129000 1720000 1 180 $X=11104000 $Y=1720000
X953 24 928 inv02 $T=11112000 3112000 0 0 $X=11112000 $Y=3112000
X954 24 929 inv02 $T=11120000 792000 0 0 $X=11120000 $Y=792000
X955 24 930 inv02 $T=11145000 1488000 1 180 $X=11120000 $Y=1488000
X956 24 931 inv02 $T=11145000 13088000 1 180 $X=11120000 $Y=13088000
X957 24 932 inv02 $T=11136000 13320000 0 0 $X=11136000 $Y=13320000
X958 24 933 inv02 $T=11169000 3112000 1 180 $X=11144000 $Y=3112000
X959 24 934 inv02 $T=11160000 560000 0 0 $X=11160000 $Y=560000
X960 24 935 inv02 $T=11176000 11464000 0 0 $X=11176000 $Y=11464000
X961 24 936 inv02 $T=11192000 560000 0 0 $X=11192000 $Y=560000
X962 24 937 inv02 $T=11200000 1720000 0 0 $X=11200000 $Y=1720000
X963 24 938 inv02 $T=11249000 6128000 1 180 $X=11224000 $Y=6128000
X964 24 939 inv02 $T=11232000 1720000 0 0 $X=11232000 $Y=1720000
X965 24 940 inv02 $T=11257000 13088000 1 180 $X=11232000 $Y=13088000
X966 24 941 inv02 $T=11264000 1720000 0 0 $X=11264000 $Y=1720000
X967 24 942 inv02 $T=11264000 9840000 0 0 $X=11264000 $Y=9840000
X968 24 943 inv02 $T=11264000 13088000 0 0 $X=11264000 $Y=13088000
X969 24 944 inv02 $T=11297000 1024000 1 180 $X=11272000 $Y=1024000
X970 24 945 inv02 $T=11280000 13320000 0 0 $X=11280000 $Y=13320000
X971 24 946 inv02 $T=11321000 1488000 1 180 $X=11296000 $Y=1488000
X972 24 947 inv02 $T=11321000 9840000 1 180 $X=11296000 $Y=9840000
X973 24 948 inv02 $T=11328000 4040000 0 0 $X=11328000 $Y=4040000
X974 24 949 inv02 $T=11328000 6592000 0 0 $X=11328000 $Y=6592000
X975 24 950 inv02 $T=11344000 9608000 0 0 $X=11344000 $Y=9608000
X976 24 951 inv02 $T=11360000 12624000 0 0 $X=11360000 $Y=12624000
X977 24 952 inv02 $T=11472000 13320000 0 0 $X=11472000 $Y=13320000
X978 24 953 inv02 $T=11528000 2648000 0 0 $X=11528000 $Y=2648000
X979 24 954 inv02 $T=11536000 1024000 0 0 $X=11536000 $Y=1024000
X980 24 955 inv02 $T=11561000 5432000 1 180 $X=11536000 $Y=5432000
X981 24 956 inv02 $T=11544000 2416000 0 0 $X=11544000 $Y=2416000
X982 24 957 inv02 $T=11577000 10072000 1 180 $X=11552000 $Y=10072000
X983 24 958 inv02 $T=11568000 1024000 0 0 $X=11568000 $Y=1024000
X984 24 959 inv02 $T=11584000 10072000 0 0 $X=11584000 $Y=10072000
X985 24 960 inv02 $T=11600000 1024000 0 0 $X=11600000 $Y=1024000
X986 24 961 inv02 $T=11616000 10072000 0 0 $X=11616000 $Y=10072000
X987 24 962 inv02 $T=11648000 5896000 0 0 $X=11648000 $Y=5896000
X988 24 963 inv02 $T=11656000 10768000 0 0 $X=11656000 $Y=10768000
X989 24 964 inv02 $T=11680000 2648000 0 0 $X=11680000 $Y=2648000
X990 24 965 inv02 $T=11680000 5896000 0 0 $X=11680000 $Y=5896000
X991 24 966 inv02 $T=11688000 10768000 0 0 $X=11688000 $Y=10768000
X992 24 967 inv02 $T=11728000 2880000 0 0 $X=11728000 $Y=2880000
X993 24 968 inv02 $T=11728000 12856000 0 0 $X=11728000 $Y=12856000
X994 24 969 inv02 $T=11744000 1488000 0 0 $X=11744000 $Y=1488000
X995 24 970 inv02 $T=11760000 7752000 0 0 $X=11760000 $Y=7752000
X996 24 971 inv02 $T=11776000 1488000 0 0 $X=11776000 $Y=1488000
X997 24 972 inv02 $T=11809000 7056000 1 180 $X=11784000 $Y=7056000
X998 24 973 inv02 $T=11817000 1024000 1 180 $X=11792000 $Y=1024000
X999 24 974 inv02 $T=11816000 5432000 0 0 $X=11816000 $Y=5432000
X1000 24 975 inv02 $T=11824000 1024000 0 0 $X=11824000 $Y=1024000
X1001 24 976 inv02 $T=11865000 560000 1 180 $X=11840000 $Y=560000
X1002 24 977 inv02 $T=11856000 1024000 0 0 $X=11856000 $Y=1024000
X1003 24 978 inv02 $T=11872000 560000 0 0 $X=11872000 $Y=560000
X1004 24 979 inv02 $T=11905000 1256000 1 180 $X=11880000 $Y=1256000
X1005 24 980 inv02 $T=11880000 4504000 0 0 $X=11880000 $Y=4504000
X1006 24 981 inv02 $T=11904000 560000 0 0 $X=11904000 $Y=560000
X1007 24 982 inv02 $T=11912000 1256000 0 0 $X=11912000 $Y=1256000
X1008 24 983 inv02 $T=11952000 1024000 0 0 $X=11952000 $Y=1024000
X1009 24 984 inv02 $T=11952000 1488000 0 0 $X=11952000 $Y=1488000
X1010 24 985 inv02 $T=11960000 7056000 0 0 $X=11960000 $Y=7056000
X1011 24 986 inv02 $T=11992000 13088000 0 0 $X=11992000 $Y=13088000
X1012 24 987 inv02 $T=12000000 11696000 0 0 $X=12000000 $Y=11696000
X1013 24 988 inv02 $T=12080000 560000 0 0 $X=12080000 $Y=560000
X1014 24 989 inv02 $T=12105000 1024000 1 180 $X=12080000 $Y=1024000
X1015 24 990 inv02 $T=12112000 560000 0 0 $X=12112000 $Y=560000
X1016 24 991 inv02 $T=12112000 1024000 0 0 $X=12112000 $Y=1024000
X1017 24 992 inv02 $T=12169000 560000 1 180 $X=12144000 $Y=560000
X1018 24 993 inv02 $T=12176000 560000 0 0 $X=12176000 $Y=560000
X1019 24 994 inv02 $T=12208000 560000 0 0 $X=12208000 $Y=560000
X1020 24 995 inv02 $T=12329000 560000 1 180 $X=12304000 $Y=560000
X1021 24 996 inv02 $T=12417000 560000 1 180 $X=12392000 $Y=560000
X1022 24 997 inv02 $T=12416000 1720000 0 0 $X=12416000 $Y=1720000
X1023 24 998 inv02 $T=12456000 1024000 0 0 $X=12456000 $Y=1024000
X1024 24 999 mux21_ni $T=152000 3344000 0 0 $X=152000 $Y=3344000
X1025 24 1000 mux21_ni $T=152000 3576000 0 0 $X=152000 $Y=3576000
X1026 24 1001 mux21_ni $T=152000 4040000 0 0 $X=152000 $Y=4040000
X1027 24 1002 mux21_ni $T=212000 4504000 1 180 $X=152000 $Y=4504000
X1028 24 1003 mux21_ni $T=152000 10304000 0 0 $X=152000 $Y=10304000
X1029 24 1004 mux21_ni $T=152000 10768000 0 0 $X=152000 $Y=10768000
X1030 24 1005 mux21_ni $T=152000 11232000 0 0 $X=152000 $Y=11232000
X1031 24 1006 mux21_ni $T=212000 11928000 1 180 $X=152000 $Y=11928000
X1032 24 1007 mux21_ni $T=152000 12624000 0 0 $X=152000 $Y=12624000
X1033 24 1008 mux21_ni $T=212000 13088000 1 180 $X=152000 $Y=13088000
X1034 24 1009 mux21_ni $T=232000 9840000 0 0 $X=232000 $Y=9840000
X1035 24 1010 mux21_ni $T=340000 2648000 1 180 $X=280000 $Y=2648000
X1036 24 1011 mux21_ni $T=280000 3576000 0 0 $X=280000 $Y=3576000
X1037 24 1012 mux21_ni $T=372000 96000 1 180 $X=312000 $Y=96000
X1038 24 1013 mux21_ni $T=372000 560000 1 180 $X=312000 $Y=560000
X1039 24 1014 mux21_ni $T=372000 792000 1 180 $X=312000 $Y=792000
X1040 24 1015 mux21_ni $T=372000 1024000 1 180 $X=312000 $Y=1024000
X1041 24 1016 mux21_ni $T=372000 1256000 1 180 $X=312000 $Y=1256000
X1042 24 1017 mux21_ni $T=372000 1488000 1 180 $X=312000 $Y=1488000
X1043 24 1018 mux21_ni $T=388000 328000 1 180 $X=328000 $Y=328000
X1044 24 1019 mux21_ni $T=336000 4040000 0 0 $X=336000 $Y=4040000
X1045 24 1020 mux21_ni $T=404000 1720000 1 180 $X=344000 $Y=1720000
X1046 24 1021 mux21_ni $T=344000 1952000 0 0 $X=344000 $Y=1952000
X1047 24 1022 mux21_ni $T=368000 4272000 0 0 $X=368000 $Y=4272000
X1048 24 1023 mux21_ni $T=428000 6360000 1 180 $X=368000 $Y=6360000
X1049 24 1024 mux21_ni $T=376000 96000 0 0 $X=376000 $Y=96000
X1050 24 1025 mux21_ni $T=436000 560000 1 180 $X=376000 $Y=560000
X1051 24 1026 mux21_ni $T=436000 1024000 1 180 $X=376000 $Y=1024000
X1052 24 1027 mux21_ni $T=436000 1488000 1 180 $X=376000 $Y=1488000
X1053 24 1028 mux21_ni $T=376000 3344000 0 0 $X=376000 $Y=3344000
X1054 24 1029 mux21_ni $T=376000 3576000 0 0 $X=376000 $Y=3576000
X1055 24 1030 mux21_ni $T=436000 8680000 1 180 $X=376000 $Y=8680000
X1056 24 1031 mux21_ni $T=460000 4736000 1 180 $X=400000 $Y=4736000
X1057 24 1032 mux21_ni $T=460000 5432000 1 180 $X=400000 $Y=5432000
X1058 24 1033 mux21_ni $T=460000 5664000 1 180 $X=400000 $Y=5664000
X1059 24 1034 mux21_ni $T=460000 7056000 1 180 $X=400000 $Y=7056000
X1060 24 1035 mux21_ni $T=460000 7520000 1 180 $X=400000 $Y=7520000
X1061 24 1036 mux21_ni $T=400000 8216000 0 0 $X=400000 $Y=8216000
X1062 24 1037 mux21_ni $T=468000 1720000 1 180 $X=408000 $Y=1720000
X1063 24 1038 mux21_ni $T=432000 2184000 0 0 $X=432000 $Y=2184000
X1064 24 1039 mux21_ni $T=440000 96000 0 0 $X=440000 $Y=96000
X1065 24 1040 mux21_ni $T=500000 560000 1 180 $X=440000 $Y=560000
X1066 24 1041 mux21_ni $T=500000 1024000 1 180 $X=440000 $Y=1024000
X1067 24 1042 mux21_ni $T=440000 1488000 0 0 $X=440000 $Y=1488000
X1068 24 1043 mux21_ni $T=500000 13320000 1 180 $X=440000 $Y=13320000
X1069 24 1044 mux21_ni $T=464000 4504000 0 0 $X=464000 $Y=4504000
X1070 24 1045 mux21_ni $T=464000 4736000 0 0 $X=464000 $Y=4736000
X1071 24 1046 mux21_ni $T=524000 5664000 1 180 $X=464000 $Y=5664000
X1072 24 1047 mux21_ni $T=532000 1720000 1 180 $X=472000 $Y=1720000
X1073 24 1048 mux21_ni $T=496000 1256000 0 0 $X=496000 $Y=1256000
X1074 24 1049 mux21_ni $T=556000 9608000 1 180 $X=496000 $Y=9608000
X1075 24 1050 mux21_ni $T=564000 96000 1 180 $X=504000 $Y=96000
X1076 24 1051 mux21_ni $T=504000 792000 0 0 $X=504000 $Y=792000
X1077 24 1052 mux21_ni $T=564000 1024000 1 180 $X=504000 $Y=1024000
X1078 24 1053 mux21_ni $T=504000 1488000 0 0 $X=504000 $Y=1488000
X1079 24 1054 mux21_ni $T=504000 2880000 0 0 $X=504000 $Y=2880000
X1080 24 1055 mux21_ni $T=504000 10304000 0 0 $X=504000 $Y=10304000
X1081 24 1056 mux21_ni $T=596000 2648000 1 180 $X=536000 $Y=2648000
X1082 24 1057 mux21_ni $T=612000 5200000 1 180 $X=552000 $Y=5200000
X1083 24 1058 mux21_ni $T=560000 12624000 0 0 $X=560000 $Y=12624000
X1084 24 1059 mux21_ni $T=568000 2880000 0 0 $X=568000 $Y=2880000
X1085 24 1060 mux21_ni $T=568000 13320000 0 0 $X=568000 $Y=13320000
X1086 24 1061 mux21_ni $T=644000 2416000 1 180 $X=584000 $Y=2416000
X1087 24 1062 mux21_ni $T=584000 7288000 0 0 $X=584000 $Y=7288000
X1088 24 1063 mux21_ni $T=600000 2648000 0 0 $X=600000 $Y=2648000
X1089 24 1064 mux21_ni $T=608000 3344000 0 0 $X=608000 $Y=3344000
X1090 24 1065 mux21_ni $T=684000 9144000 1 180 $X=624000 $Y=9144000
X1091 24 1066 mux21_ni $T=632000 3808000 0 0 $X=632000 $Y=3808000
X1092 24 1067 mux21_ni $T=640000 5896000 0 0 $X=640000 $Y=5896000
X1093 24 1068 mux21_ni $T=672000 3344000 0 0 $X=672000 $Y=3344000
X1094 24 1069 mux21_ni $T=680000 5664000 0 0 $X=680000 $Y=5664000
X1095 24 1070 mux21_ni $T=748000 9144000 1 180 $X=688000 $Y=9144000
X1096 24 1071 mux21_ni $T=764000 11464000 1 180 $X=704000 $Y=11464000
X1097 24 1072 mux21_ni $T=712000 10072000 0 0 $X=712000 $Y=10072000
X1098 24 1073 mux21_ni $T=720000 1952000 0 0 $X=720000 $Y=1952000
X1099 24 1074 mux21_ni $T=720000 7984000 0 0 $X=720000 $Y=7984000
X1100 24 1075 mux21_ni $T=736000 6360000 0 0 $X=736000 $Y=6360000
X1101 24 1076 mux21_ni $T=804000 1720000 1 180 $X=744000 $Y=1720000
X1102 24 1077 mux21_ni $T=744000 2184000 0 0 $X=744000 $Y=2184000
X1103 24 1078 mux21_ni $T=744000 4504000 0 0 $X=744000 $Y=4504000
X1104 24 1079 mux21_ni $T=844000 560000 1 180 $X=784000 $Y=560000
X1105 24 1080 mux21_ni $T=844000 1952000 1 180 $X=784000 $Y=1952000
X1106 24 1081 mux21_ni $T=792000 96000 0 0 $X=792000 $Y=96000
X1107 24 1082 mux21_ni $T=852000 7752000 1 180 $X=792000 $Y=7752000
X1108 24 1083 mux21_ni $T=816000 4736000 0 0 $X=816000 $Y=4736000
X1109 24 1084 mux21_ni $T=884000 328000 1 180 $X=824000 $Y=328000
X1110 24 1085 mux21_ni $T=884000 2648000 1 180 $X=824000 $Y=2648000
X1111 24 1086 mux21_ni $T=884000 9608000 1 180 $X=824000 $Y=9608000
X1112 24 1087 mux21_ni $T=908000 560000 1 180 $X=848000 $Y=560000
X1113 24 1088 mux21_ni $T=848000 792000 0 0 $X=848000 $Y=792000
X1114 24 1089 mux21_ni $T=848000 1024000 0 0 $X=848000 $Y=1024000
X1115 24 1090 mux21_ni $T=908000 1952000 1 180 $X=848000 $Y=1952000
X1116 24 1091 mux21_ni $T=856000 1488000 0 0 $X=856000 $Y=1488000
X1117 24 1092 mux21_ni $T=888000 6360000 0 0 $X=888000 $Y=6360000
X1118 24 1093 mux21_ni $T=964000 7752000 1 180 $X=904000 $Y=7752000
X1119 24 1094 mux21_ni $T=912000 2416000 0 0 $X=912000 $Y=2416000
X1120 24 1095 mux21_ni $T=912000 5432000 0 0 $X=912000 $Y=5432000
X1121 24 1096 mux21_ni $T=920000 1488000 0 0 $X=920000 $Y=1488000
X1122 24 1097 mux21_ni $T=920000 4968000 0 0 $X=920000 $Y=4968000
X1123 24 1098 mux21_ni $T=980000 11696000 1 180 $X=920000 $Y=11696000
X1124 24 1099 mux21_ni $T=928000 13552000 0 0 $X=928000 $Y=13552000
X1125 24 1100 mux21_ni $T=1004000 12392000 1 180 $X=944000 $Y=12392000
X1126 24 1101 mux21_ni $T=1012000 7288000 1 180 $X=952000 $Y=7288000
X1127 24 1102 mux21_ni $T=1028000 1720000 1 180 $X=968000 $Y=1720000
X1128 24 1103 mux21_ni $T=968000 10304000 0 0 $X=968000 $Y=10304000
X1129 24 1104 mux21_ni $T=976000 792000 0 0 $X=976000 $Y=792000
X1130 24 1105 mux21_ni $T=976000 2416000 0 0 $X=976000 $Y=2416000
X1131 24 1106 mux21_ni $T=984000 1488000 0 0 $X=984000 $Y=1488000
X1132 24 1107 mux21_ni $T=984000 11232000 0 0 $X=984000 $Y=11232000
X1133 24 1108 mux21_ni $T=984000 13088000 0 0 $X=984000 $Y=13088000
X1134 24 1109 mux21_ni $T=1092000 1720000 1 180 $X=1032000 $Y=1720000
X1135 24 1110 mux21_ni $T=1040000 2416000 0 0 $X=1040000 $Y=2416000
X1136 24 1111 mux21_ni $T=1040000 12160000 0 0 $X=1040000 $Y=12160000
X1137 24 1112 mux21_ni $T=1048000 1488000 0 0 $X=1048000 $Y=1488000
X1138 24 1113 mux21_ni $T=1048000 5664000 0 0 $X=1048000 $Y=5664000
X1139 24 1114 mux21_ni $T=1064000 11696000 0 0 $X=1064000 $Y=11696000
X1140 24 1115 mux21_ni $T=1072000 1024000 0 0 $X=1072000 $Y=1024000
X1141 24 1116 mux21_ni $T=1132000 4040000 1 180 $X=1072000 $Y=4040000
X1142 24 1117 mux21_ni $T=1140000 328000 1 180 $X=1080000 $Y=328000
X1143 24 1118 mux21_ni $T=1148000 3344000 1 180 $X=1088000 $Y=3344000
X1144 24 1119 mux21_ni $T=1188000 1720000 1 180 $X=1128000 $Y=1720000
X1145 24 1120 mux21_ni $T=1128000 12624000 0 0 $X=1128000 $Y=12624000
X1146 24 1121 mux21_ni $T=1136000 1024000 0 0 $X=1136000 $Y=1024000
X1147 24 1122 mux21_ni $T=1136000 4040000 0 0 $X=1136000 $Y=4040000
X1148 24 1123 mux21_ni $T=1212000 3576000 1 180 $X=1152000 $Y=3576000
X1149 24 1124 mux21_ni $T=1168000 11928000 0 0 $X=1168000 $Y=11928000
X1150 24 1125 mux21_ni $T=1252000 1720000 1 180 $X=1192000 $Y=1720000
X1151 24 1126 mux21_ni $T=1252000 3808000 1 180 $X=1192000 $Y=3808000
X1152 24 1127 mux21_ni $T=1192000 6360000 0 0 $X=1192000 $Y=6360000
X1153 24 1128 mux21_ni $T=1260000 560000 1 180 $X=1200000 $Y=560000
X1154 24 1129 mux21_ni $T=1284000 13320000 1 180 $X=1224000 $Y=13320000
X1155 24 1130 mux21_ni $T=1232000 11464000 0 0 $X=1232000 $Y=11464000
X1156 24 1131 mux21_ni $T=1248000 10536000 0 0 $X=1248000 $Y=10536000
X1157 24 1132 mux21_ni $T=1256000 1720000 0 0 $X=1256000 $Y=1720000
X1158 24 1133 mux21_ni $T=1316000 3808000 1 180 $X=1256000 $Y=3808000
X1159 24 1134 mux21_ni $T=1256000 4040000 0 0 $X=1256000 $Y=4040000
X1160 24 1135 mux21_ni $T=1288000 13088000 0 0 $X=1288000 $Y=13088000
X1161 24 1136 mux21_ni $T=1296000 11464000 0 0 $X=1296000 $Y=11464000
X1162 24 1137 mux21_ni $T=1380000 1720000 1 180 $X=1320000 $Y=1720000
X1163 24 1138 mux21_ni $T=1328000 10304000 0 0 $X=1328000 $Y=10304000
X1164 24 1139 mux21_ni $T=1328000 13320000 0 0 $X=1328000 $Y=13320000
X1165 24 1140 mux21_ni $T=1344000 3576000 0 0 $X=1344000 $Y=3576000
X1166 24 1141 mux21_ni $T=1344000 5200000 0 0 $X=1344000 $Y=5200000
X1167 24 1142 mux21_ni $T=1352000 12856000 0 0 $X=1352000 $Y=12856000
X1168 24 1143 mux21_ni $T=1376000 11232000 0 0 $X=1376000 $Y=11232000
X1169 24 1144 mux21_ni $T=1476000 96000 1 180 $X=1416000 $Y=96000
X1170 24 1145 mux21_ni $T=1492000 1488000 1 180 $X=1432000 $Y=1488000
X1171 24 1146 mux21_ni $T=1432000 7056000 0 0 $X=1432000 $Y=7056000
X1172 24 1147 mux21_ni $T=1508000 3808000 1 180 $X=1448000 $Y=3808000
X1173 24 1148 mux21_ni $T=1516000 6824000 1 180 $X=1456000 $Y=6824000
X1174 24 1149 mux21_ni $T=1524000 1256000 1 180 $X=1464000 $Y=1256000
X1175 24 1150 mux21_ni $T=1540000 96000 1 180 $X=1480000 $Y=96000
X1176 24 1151 mux21_ni $T=1548000 560000 1 180 $X=1488000 $Y=560000
X1177 24 1152 mux21_ni $T=1496000 2184000 0 0 $X=1496000 $Y=2184000
X1178 24 1153 mux21_ni $T=1504000 6360000 0 0 $X=1504000 $Y=6360000
X1179 24 1154 mux21_ni $T=1512000 3808000 0 0 $X=1512000 $Y=3808000
X1180 24 1155 mux21_ni $T=1520000 6824000 0 0 $X=1520000 $Y=6824000
X1181 24 1156 mux21_ni $T=1520000 12392000 0 0 $X=1520000 $Y=12392000
X1182 24 1157 mux21_ni $T=1588000 328000 1 180 $X=1528000 $Y=328000
X1183 24 1158 mux21_ni $T=1528000 1256000 0 0 $X=1528000 $Y=1256000
X1184 24 1159 mux21_ni $T=1604000 96000 1 180 $X=1544000 $Y=96000
X1185 24 1160 mux21_ni $T=1612000 560000 1 180 $X=1552000 $Y=560000
X1186 24 1161 mux21_ni $T=1612000 1024000 1 180 $X=1552000 $Y=1024000
X1187 24 1162 mux21_ni $T=1552000 8216000 0 0 $X=1552000 $Y=8216000
X1188 24 1163 mux21_ni $T=1568000 7288000 0 0 $X=1568000 $Y=7288000
X1189 24 1164 mux21_ni $T=1568000 7984000 0 0 $X=1568000 $Y=7984000
X1190 24 1165 mux21_ni $T=1576000 3808000 0 0 $X=1576000 $Y=3808000
X1191 24 1166 mux21_ni $T=1584000 3344000 0 0 $X=1584000 $Y=3344000
X1192 24 1167 mux21_ni $T=1584000 6824000 0 0 $X=1584000 $Y=6824000
X1193 24 1168 mux21_ni $T=1592000 328000 0 0 $X=1592000 $Y=328000
X1194 24 1169 mux21_ni $T=1592000 6592000 0 0 $X=1592000 $Y=6592000
X1195 24 1170 mux21_ni $T=1600000 3576000 0 0 $X=1600000 $Y=3576000
X1196 24 1171 mux21_ni $T=1608000 5896000 0 0 $X=1608000 $Y=5896000
X1197 24 1172 mux21_ni $T=1608000 7752000 0 0 $X=1608000 $Y=7752000
X1198 24 1173 mux21_ni $T=1616000 1024000 0 0 $X=1616000 $Y=1024000
X1199 24 1174 mux21_ni $T=1624000 8448000 0 0 $X=1624000 $Y=8448000
X1200 24 1175 mux21_ni $T=1708000 6824000 1 180 $X=1648000 $Y=6824000
X1201 24 1176 mux21_ni $T=1716000 328000 1 180 $X=1656000 $Y=328000
X1202 24 1177 mux21_ni $T=1656000 5664000 0 0 $X=1656000 $Y=5664000
X1203 24 1178 mux21_ni $T=1740000 11000000 1 180 $X=1680000 $Y=11000000
X1204 24 1179 mux21_ni $T=1688000 6128000 0 0 $X=1688000 $Y=6128000
X1205 24 1180 mux21_ni $T=1688000 7056000 0 0 $X=1688000 $Y=7056000
X1206 24 1181 mux21_ni $T=1688000 7520000 0 0 $X=1688000 $Y=7520000
X1207 24 1182 mux21_ni $T=1688000 11232000 0 0 $X=1688000 $Y=11232000
X1208 24 1183 mux21_ni $T=1756000 792000 1 180 $X=1696000 $Y=792000
X1209 24 1184 mux21_ni $T=1704000 5432000 0 0 $X=1704000 $Y=5432000
X1210 24 1185 mux21_ni $T=1704000 10304000 0 0 $X=1704000 $Y=10304000
X1211 24 1186 mux21_ni $T=1736000 6824000 0 0 $X=1736000 $Y=6824000
X1212 24 1187 mux21_ni $T=1804000 1952000 1 180 $X=1744000 $Y=1952000
X1213 24 1188 mux21_ni $T=1752000 1488000 0 0 $X=1752000 $Y=1488000
X1214 24 1189 mux21_ni $T=1752000 10536000 0 0 $X=1752000 $Y=10536000
X1215 24 1190 mux21_ni $T=1820000 792000 1 180 $X=1760000 $Y=792000
X1216 24 1191 mux21_ni $T=1820000 13552000 1 180 $X=1760000 $Y=13552000
X1217 24 1192 mux21_ni $T=1828000 96000 1 180 $X=1768000 $Y=96000
X1218 24 1193 mux21_ni $T=1808000 560000 0 0 $X=1808000 $Y=560000
X1219 24 1194 mux21_ni $T=1816000 1488000 0 0 $X=1816000 $Y=1488000
X1220 24 1195 mux21_ni $T=1816000 4504000 0 0 $X=1816000 $Y=4504000
X1221 24 1196 mux21_ni $T=1876000 10072000 1 180 $X=1816000 $Y=10072000
X1222 24 1197 mux21_ni $T=1824000 13552000 0 0 $X=1824000 $Y=13552000
X1223 24 1198 mux21_ni $T=1892000 4272000 1 180 $X=1832000 $Y=4272000
X1224 24 1199 mux21_ni $T=1832000 4968000 0 0 $X=1832000 $Y=4968000
X1225 24 1200 mux21_ni $T=1840000 1024000 0 0 $X=1840000 $Y=1024000
X1226 24 1201 mux21_ni $T=1856000 1952000 0 0 $X=1856000 $Y=1952000
X1227 24 1202 mux21_ni $T=1864000 3344000 0 0 $X=1864000 $Y=3344000
X1228 24 1203 mux21_ni $T=1924000 13088000 1 180 $X=1864000 $Y=13088000
X1229 24 1204 mux21_ni $T=1880000 13320000 0 0 $X=1880000 $Y=13320000
X1230 24 1205 mux21_ni $T=1888000 8912000 0 0 $X=1888000 $Y=8912000
X1231 24 1206 mux21_ni $T=1904000 1024000 0 0 $X=1904000 $Y=1024000
X1232 24 1207 mux21_ni $T=1904000 9144000 0 0 $X=1904000 $Y=9144000
X1233 24 1208 mux21_ni $T=1912000 8216000 0 0 $X=1912000 $Y=8216000
X1234 24 1209 mux21_ni $T=1928000 8448000 0 0 $X=1928000 $Y=8448000
X1235 24 1210 mux21_ni $T=1928000 8680000 0 0 $X=1928000 $Y=8680000
X1236 24 1211 mux21_ni $T=2020000 3112000 1 180 $X=1960000 $Y=3112000
X1237 24 1212 mux21_ni $T=1960000 9608000 0 0 $X=1960000 $Y=9608000
X1238 24 1213 mux21_ni $T=2052000 96000 1 180 $X=1992000 $Y=96000
X1239 24 1214 mux21_ni $T=2060000 328000 1 180 $X=2000000 $Y=328000
X1240 24 1215 mux21_ni $T=2016000 1256000 0 0 $X=2016000 $Y=1256000
X1241 24 1216 mux21_ni $T=2092000 1720000 1 180 $X=2032000 $Y=1720000
X1242 24 1217 mux21_ni $T=2092000 12392000 1 180 $X=2032000 $Y=12392000
X1243 24 1218 mux21_ni $T=2040000 1024000 0 0 $X=2040000 $Y=1024000
X1244 24 1219 mux21_ni $T=2116000 96000 1 180 $X=2056000 $Y=96000
X1245 24 1220 mux21_ni $T=2124000 328000 1 180 $X=2064000 $Y=328000
X1246 24 1221 mux21_ni $T=2132000 7288000 1 180 $X=2072000 $Y=7288000
X1247 24 1222 mux21_ni $T=2080000 1952000 0 0 $X=2080000 $Y=1952000
X1248 24 1223 mux21_ni $T=2080000 2184000 0 0 $X=2080000 $Y=2184000
X1249 24 1224 mux21_ni $T=2096000 13088000 0 0 $X=2096000 $Y=13088000
X1250 24 1225 mux21_ni $T=2104000 6128000 0 0 $X=2104000 $Y=6128000
X1251 24 1226 mux21_ni $T=2136000 4968000 0 0 $X=2136000 $Y=4968000
X1252 24 1227 mux21_ni $T=2136000 6360000 0 0 $X=2136000 $Y=6360000
X1253 24 1228 mux21_ni $T=2136000 7288000 0 0 $X=2136000 $Y=7288000
X1254 24 1229 mux21_ni $T=2144000 1256000 0 0 $X=2144000 $Y=1256000
X1255 24 1230 mux21_ni $T=2168000 4504000 0 0 $X=2168000 $Y=4504000
X1256 24 1231 mux21_ni $T=2176000 6592000 0 0 $X=2176000 $Y=6592000
X1257 24 1232 mux21_ni $T=2184000 3808000 0 0 $X=2184000 $Y=3808000
X1258 24 1233 mux21_ni $T=2192000 8912000 0 0 $X=2192000 $Y=8912000
X1259 24 1234 mux21_ni $T=2208000 1256000 0 0 $X=2208000 $Y=1256000
X1260 24 1235 mux21_ni $T=2208000 4272000 0 0 $X=2208000 $Y=4272000
X1261 24 1236 mux21_ni $T=2216000 7056000 0 0 $X=2216000 $Y=7056000
X1262 24 1237 mux21_ni $T=2224000 7752000 0 0 $X=2224000 $Y=7752000
X1263 24 1238 mux21_ni $T=2232000 2648000 0 0 $X=2232000 $Y=2648000
X1264 24 1239 mux21_ni $T=2288000 792000 0 0 $X=2288000 $Y=792000
X1265 24 1240 mux21_ni $T=2288000 7752000 0 0 $X=2288000 $Y=7752000
X1266 24 1241 mux21_ni $T=2288000 11000000 0 0 $X=2288000 $Y=11000000
X1267 24 1242 mux21_ni $T=2312000 5432000 0 0 $X=2312000 $Y=5432000
X1268 24 1243 mux21_ni $T=2336000 560000 0 0 $X=2336000 $Y=560000
X1269 24 1244 mux21_ni $T=2352000 9144000 0 0 $X=2352000 $Y=9144000
X1270 24 1245 mux21_ni $T=2420000 3344000 1 180 $X=2360000 $Y=3344000
X1271 24 1246 mux21_ni $T=2444000 96000 1 180 $X=2384000 $Y=96000
X1272 24 1247 mux21_ni $T=2460000 5664000 1 180 $X=2400000 $Y=5664000
X1273 24 1248 mux21_ni $T=2468000 328000 1 180 $X=2408000 $Y=328000
X1274 24 1249 mux21_ni $T=2408000 4040000 0 0 $X=2408000 $Y=4040000
X1275 24 1250 mux21_ni $T=2408000 6128000 0 0 $X=2408000 $Y=6128000
X1276 24 1251 mux21_ni $T=2468000 13320000 1 180 $X=2408000 $Y=13320000
X1277 24 1252 mux21_ni $T=2432000 1256000 0 0 $X=2432000 $Y=1256000
X1278 24 1253 mux21_ni $T=2432000 10536000 0 0 $X=2432000 $Y=10536000
X1279 24 1254 mux21_ni $T=2508000 96000 1 180 $X=2448000 $Y=96000
X1280 24 1255 mux21_ni $T=2516000 4736000 1 180 $X=2456000 $Y=4736000
X1281 24 1256 mux21_ni $T=2472000 328000 0 0 $X=2472000 $Y=328000
X1282 24 1257 mux21_ni $T=2496000 1256000 0 0 $X=2496000 $Y=1256000
X1283 24 1258 mux21_ni $T=2572000 96000 1 180 $X=2512000 $Y=96000
X1284 24 1259 mux21_ni $T=2512000 1024000 0 0 $X=2512000 $Y=1024000
X1285 24 1260 mux21_ni $T=2528000 7056000 0 0 $X=2528000 $Y=7056000
X1286 24 1261 mux21_ni $T=2596000 328000 1 180 $X=2536000 $Y=328000
X1287 24 1262 mux21_ni $T=2544000 1720000 0 0 $X=2544000 $Y=1720000
X1288 24 1263 mux21_ni $T=2604000 12624000 1 180 $X=2544000 $Y=12624000
X1289 24 1264 mux21_ni $T=2604000 12856000 1 180 $X=2544000 $Y=12856000
X1290 24 1265 mux21_ni $T=2620000 560000 1 180 $X=2560000 $Y=560000
X1291 24 1266 mux21_ni $T=2568000 4272000 0 0 $X=2568000 $Y=4272000
X1292 24 1267 mux21_ni $T=2636000 96000 1 180 $X=2576000 $Y=96000
X1293 24 1268 mux21_ni $T=2584000 5200000 0 0 $X=2584000 $Y=5200000
X1294 24 1269 mux21_ni $T=2592000 7752000 0 0 $X=2592000 $Y=7752000
X1295 24 1270 mux21_ni $T=2600000 328000 0 0 $X=2600000 $Y=328000
X1296 24 1271 mux21_ni $T=2624000 5432000 0 0 $X=2624000 $Y=5432000
X1297 24 1272 mux21_ni $T=2648000 12160000 0 0 $X=2648000 $Y=12160000
X1298 24 1273 mux21_ni $T=2656000 3112000 0 0 $X=2656000 $Y=3112000
X1299 24 1274 mux21_ni $T=2656000 8216000 0 0 $X=2656000 $Y=8216000
X1300 24 1275 mux21_ni $T=2672000 792000 0 0 $X=2672000 $Y=792000
X1301 24 1276 mux21_ni $T=2740000 12856000 1 180 $X=2680000 $Y=12856000
X1302 24 1277 mux21_ni $T=2764000 1952000 1 180 $X=2704000 $Y=1952000
X1303 24 1278 mux21_ni $T=2712000 4040000 0 0 $X=2712000 $Y=4040000
X1304 24 1279 mux21_ni $T=2728000 10304000 0 0 $X=2728000 $Y=10304000
X1305 24 1280 mux21_ni $T=2736000 792000 0 0 $X=2736000 $Y=792000
X1306 24 1281 mux21_ni $T=2796000 1024000 1 180 $X=2736000 $Y=1024000
X1307 24 1282 mux21_ni $T=2736000 3576000 0 0 $X=2736000 $Y=3576000
X1308 24 1283 mux21_ni $T=2752000 3344000 0 0 $X=2752000 $Y=3344000
X1309 24 1284 mux21_ni $T=2752000 6824000 0 0 $X=2752000 $Y=6824000
X1310 24 1285 mux21_ni $T=2828000 13320000 1 180 $X=2768000 $Y=13320000
X1311 24 1286 mux21_ni $T=2844000 1256000 1 180 $X=2784000 $Y=1256000
X1312 24 1287 mux21_ni $T=2844000 1488000 1 180 $X=2784000 $Y=1488000
X1313 24 1288 mux21_ni $T=2792000 3808000 0 0 $X=2792000 $Y=3808000
X1314 24 1289 mux21_ni $T=2908000 2184000 1 180 $X=2848000 $Y=2184000
X1315 24 1290 mux21_ni $T=2924000 96000 1 180 $X=2864000 $Y=96000
X1316 24 1291 mux21_ni $T=2924000 4736000 1 180 $X=2864000 $Y=4736000
X1317 24 1292 mux21_ni $T=2924000 8912000 1 180 $X=2864000 $Y=8912000
X1318 24 1293 mux21_ni $T=2872000 4272000 0 0 $X=2872000 $Y=4272000
X1319 24 1294 mux21_ni $T=2932000 4504000 1 180 $X=2872000 $Y=4504000
X1320 24 1295 mux21_ni $T=2872000 5896000 0 0 $X=2872000 $Y=5896000
X1321 24 1296 mux21_ni $T=2872000 13552000 0 0 $X=2872000 $Y=13552000
X1322 24 1297 mux21_ni $T=2888000 7288000 0 0 $X=2888000 $Y=7288000
X1323 24 1298 mux21_ni $T=2956000 9144000 1 180 $X=2896000 $Y=9144000
X1324 24 1299 mux21_ni $T=2904000 10768000 0 0 $X=2904000 $Y=10768000
X1325 24 1300 mux21_ni $T=2928000 13088000 0 0 $X=2928000 $Y=13088000
X1326 24 1301 mux21_ni $T=2928000 13320000 0 0 $X=2928000 $Y=13320000
X1327 24 1302 mux21_ni $T=2936000 5896000 0 0 $X=2936000 $Y=5896000
X1328 24 1303 mux21_ni $T=3036000 1952000 1 180 $X=2976000 $Y=1952000
X1329 24 1304 mux21_ni $T=2976000 2184000 0 0 $X=2976000 $Y=2184000
X1330 24 1305 mux21_ni $T=2984000 9840000 0 0 $X=2984000 $Y=9840000
X1331 24 1306 mux21_ni $T=2992000 4504000 0 0 $X=2992000 $Y=4504000
X1332 24 1307 mux21_ni $T=2992000 4736000 0 0 $X=2992000 $Y=4736000
X1333 24 1308 mux21_ni $T=3000000 3112000 0 0 $X=3000000 $Y=3112000
X1334 24 1309 mux21_ni $T=3008000 12856000 0 0 $X=3008000 $Y=12856000
X1335 24 1310 mux21_ni $T=3084000 12392000 1 180 $X=3024000 $Y=12392000
X1336 24 1311 mux21_ni $T=3092000 6360000 1 180 $X=3032000 $Y=6360000
X1337 24 1312 mux21_ni $T=3108000 3808000 1 180 $X=3048000 $Y=3808000
X1338 24 1313 mux21_ni $T=3140000 1024000 1 180 $X=3080000 $Y=1024000
X1339 24 1314 mux21_ni $T=3140000 2416000 1 180 $X=3080000 $Y=2416000
X1340 24 1315 mux21_ni $T=3088000 3344000 0 0 $X=3088000 $Y=3344000
X1341 24 1316 mux21_ni $T=3088000 7752000 0 0 $X=3088000 $Y=7752000
X1342 24 1317 mux21_ni $T=3088000 9376000 0 0 $X=3088000 $Y=9376000
X1343 24 1318 mux21_ni $T=3096000 3576000 0 0 $X=3096000 $Y=3576000
X1344 24 1319 mux21_ni $T=3164000 1952000 1 180 $X=3104000 $Y=1952000
X1345 24 1320 mux21_ni $T=3112000 5200000 0 0 $X=3112000 $Y=5200000
X1346 24 1321 mux21_ni $T=3120000 2880000 0 0 $X=3120000 $Y=2880000
X1347 24 1322 mux21_ni $T=3120000 5432000 0 0 $X=3120000 $Y=5432000
X1348 24 1323 mux21_ni $T=3128000 2648000 0 0 $X=3128000 $Y=2648000
X1349 24 1324 mux21_ni $T=3128000 6360000 0 0 $X=3128000 $Y=6360000
X1350 24 1325 mux21_ni $T=3128000 10304000 0 0 $X=3128000 $Y=10304000
X1351 24 1326 mux21_ni $T=3136000 560000 0 0 $X=3136000 $Y=560000
X1352 24 1327 mux21_ni $T=3144000 4968000 0 0 $X=3144000 $Y=4968000
X1353 24 1328 mux21_ni $T=3144000 10072000 0 0 $X=3144000 $Y=10072000
X1354 24 1329 mux21_ni $T=3212000 792000 1 180 $X=3152000 $Y=792000
X1355 24 1330 mux21_ni $T=3152000 4272000 0 0 $X=3152000 $Y=4272000
X1356 24 1331 mux21_ni $T=3184000 8912000 0 0 $X=3184000 $Y=8912000
X1357 24 1332 mux21_ni $T=3216000 792000 0 0 $X=3216000 $Y=792000
X1358 24 1333 mux21_ni $T=3216000 4272000 0 0 $X=3216000 $Y=4272000
X1359 24 1334 mux21_ni $T=3216000 7056000 0 0 $X=3216000 $Y=7056000
X1360 24 1335 mux21_ni $T=3216000 9608000 0 0 $X=3216000 $Y=9608000
X1361 24 1336 mux21_ni $T=3248000 5896000 0 0 $X=3248000 $Y=5896000
X1362 24 1337 mux21_ni $T=3324000 11464000 1 180 $X=3264000 $Y=11464000
X1363 24 1338 mux21_ni $T=3324000 12160000 1 180 $X=3264000 $Y=12160000
X1364 24 1339 mux21_ni $T=3280000 7056000 0 0 $X=3280000 $Y=7056000
X1365 24 1340 mux21_ni $T=3288000 6824000 0 0 $X=3288000 $Y=6824000
X1366 24 1341 mux21_ni $T=3368000 1720000 0 0 $X=3368000 $Y=1720000
X1367 24 1342 mux21_ni $T=3368000 13552000 0 0 $X=3368000 $Y=13552000
X1368 24 1343 mux21_ni $T=3392000 1024000 0 0 $X=3392000 $Y=1024000
X1369 24 1344 mux21_ni $T=3392000 2416000 0 0 $X=3392000 $Y=2416000
X1370 24 1345 mux21_ni $T=3400000 2880000 0 0 $X=3400000 $Y=2880000
X1371 24 1346 mux21_ni $T=3408000 10304000 0 0 $X=3408000 $Y=10304000
X1372 24 1347 mux21_ni $T=3416000 1952000 0 0 $X=3416000 $Y=1952000
X1373 24 1348 mux21_ni $T=3476000 3808000 1 180 $X=3416000 $Y=3808000
X1374 24 1349 mux21_ni $T=3416000 12624000 0 0 $X=3416000 $Y=12624000
X1375 24 1350 mux21_ni $T=3484000 328000 1 180 $X=3424000 $Y=328000
X1376 24 1351 mux21_ni $T=3424000 4968000 0 0 $X=3424000 $Y=4968000
X1377 24 1352 mux21_ni $T=3424000 6128000 0 0 $X=3424000 $Y=6128000
X1378 24 1353 mux21_ni $T=3432000 12856000 0 0 $X=3432000 $Y=12856000
X1379 24 1354 mux21_ni $T=3448000 2184000 0 0 $X=3448000 $Y=2184000
X1380 24 1355 mux21_ni $T=3456000 7984000 0 0 $X=3456000 $Y=7984000
X1381 24 1356 mux21_ni $T=3480000 3808000 0 0 $X=3480000 $Y=3808000
X1382 24 1357 mux21_ni $T=3528000 9144000 0 0 $X=3528000 $Y=9144000
X1383 24 1358 mux21_ni $T=3560000 8680000 0 0 $X=3560000 $Y=8680000
X1384 24 1359 mux21_ni $T=3584000 7056000 0 0 $X=3584000 $Y=7056000
X1385 24 1360 mux21_ni $T=3652000 7520000 1 180 $X=3592000 $Y=7520000
X1386 24 1361 mux21_ni $T=3680000 2648000 0 0 $X=3680000 $Y=2648000
X1387 24 1362 mux21_ni $T=3680000 9376000 0 0 $X=3680000 $Y=9376000
X1388 24 1363 mux21_ni $T=3680000 10768000 0 0 $X=3680000 $Y=10768000
X1389 24 1364 mux21_ni $T=3680000 11000000 0 0 $X=3680000 $Y=11000000
X1390 24 1365 mux21_ni $T=3688000 1488000 0 0 $X=3688000 $Y=1488000
X1391 24 1366 mux21_ni $T=3712000 7056000 0 0 $X=3712000 $Y=7056000
X1392 24 1367 mux21_ni $T=3712000 8448000 0 0 $X=3712000 $Y=8448000
X1393 24 1368 mux21_ni $T=3712000 11696000 0 0 $X=3712000 $Y=11696000
X1394 24 1369 mux21_ni $T=3720000 1952000 0 0 $X=3720000 $Y=1952000
X1395 24 1370 mux21_ni $T=3728000 2880000 0 0 $X=3728000 $Y=2880000
X1396 24 1371 mux21_ni $T=3728000 4504000 0 0 $X=3728000 $Y=4504000
X1397 24 1372 mux21_ni $T=3728000 6592000 0 0 $X=3728000 $Y=6592000
X1398 24 1373 mux21_ni $T=3744000 3112000 0 0 $X=3744000 $Y=3112000
X1399 24 1374 mux21_ni $T=3760000 4040000 0 0 $X=3760000 $Y=4040000
X1400 24 1375 mux21_ni $T=3776000 7520000 0 0 $X=3776000 $Y=7520000
X1401 24 1376 mux21_ni $T=3776000 8448000 0 0 $X=3776000 $Y=8448000
X1402 24 1377 mux21_ni $T=3784000 2416000 0 0 $X=3784000 $Y=2416000
X1403 24 1378 mux21_ni $T=3784000 3808000 0 0 $X=3784000 $Y=3808000
X1404 24 1379 mux21_ni $T=3784000 7288000 0 0 $X=3784000 $Y=7288000
X1405 24 1380 mux21_ni $T=3852000 4736000 1 180 $X=3792000 $Y=4736000
X1406 24 1381 mux21_ni $T=3816000 11928000 0 0 $X=3816000 $Y=11928000
X1407 24 1382 mux21_ni $T=3832000 328000 0 0 $X=3832000 $Y=328000
X1408 24 1383 mux21_ni $T=3840000 4968000 0 0 $X=3840000 $Y=4968000
X1409 24 1384 mux21_ni $T=3848000 6824000 0 0 $X=3848000 $Y=6824000
X1410 24 1385 mux21_ni $T=3872000 5432000 0 0 $X=3872000 $Y=5432000
X1411 24 1386 mux21_ni $T=3872000 8680000 0 0 $X=3872000 $Y=8680000
X1412 24 1387 mux21_ni $T=3896000 3344000 0 0 $X=3896000 $Y=3344000
X1413 24 1388 mux21_ni $T=3912000 4736000 0 0 $X=3912000 $Y=4736000
X1414 24 1389 mux21_ni $T=3928000 5200000 0 0 $X=3928000 $Y=5200000
X1415 24 1390 mux21_ni $T=3988000 12856000 1 180 $X=3928000 $Y=12856000
X1416 24 1391 mux21_ni $T=4004000 560000 1 180 $X=3944000 $Y=560000
X1417 24 1392 mux21_ni $T=3944000 1024000 0 0 $X=3944000 $Y=1024000
X1418 24 1393 mux21_ni $T=4036000 11232000 1 180 $X=3976000 $Y=11232000
X1419 24 1394 mux21_ni $T=4044000 10768000 1 180 $X=3984000 $Y=10768000
X1420 24 1395 mux21_ni $T=3992000 792000 0 0 $X=3992000 $Y=792000
X1421 24 1396 mux21_ni $T=3992000 10536000 0 0 $X=3992000 $Y=10536000
X1422 24 1397 mux21_ni $T=4068000 560000 1 180 $X=4008000 $Y=560000
X1423 24 1398 mux21_ni $T=4032000 6592000 0 0 $X=4032000 $Y=6592000
X1424 24 1399 mux21_ni $T=4032000 7752000 0 0 $X=4032000 $Y=7752000
X1425 24 1400 mux21_ni $T=4092000 13320000 1 180 $X=4032000 $Y=13320000
X1426 24 1401 mux21_ni $T=4040000 4272000 0 0 $X=4040000 $Y=4272000
X1427 24 1402 mux21_ni $T=4056000 10304000 0 0 $X=4056000 $Y=10304000
X1428 24 1403 mux21_ni $T=4072000 3576000 0 0 $X=4072000 $Y=3576000
X1429 24 1404 mux21_ni $T=4088000 3808000 0 0 $X=4088000 $Y=3808000
X1430 24 1405 mux21_ni $T=4088000 10768000 0 0 $X=4088000 $Y=10768000
X1431 24 1406 mux21_ni $T=4164000 1720000 1 180 $X=4104000 $Y=1720000
X1432 24 1407 mux21_ni $T=4104000 6360000 0 0 $X=4104000 $Y=6360000
X1433 24 1408 mux21_ni $T=4136000 1952000 0 0 $X=4136000 $Y=1952000
X1434 24 1409 mux21_ni $T=4136000 7520000 0 0 $X=4136000 $Y=7520000
X1435 24 1410 mux21_ni $T=4144000 2880000 0 0 $X=4144000 $Y=2880000
X1436 24 1411 mux21_ni $T=4152000 4504000 0 0 $X=4152000 $Y=4504000
X1437 24 1412 mux21_ni $T=4228000 560000 1 180 $X=4168000 $Y=560000
X1438 24 1413 mux21_ni $T=4168000 1720000 0 0 $X=4168000 $Y=1720000
X1439 24 1414 mux21_ni $T=4168000 8216000 0 0 $X=4168000 $Y=8216000
X1440 24 1415 mux21_ni $T=4176000 1256000 0 0 $X=4176000 $Y=1256000
X1441 24 1416 mux21_ni $T=4184000 1488000 0 0 $X=4184000 $Y=1488000
X1442 24 1417 mux21_ni $T=4232000 560000 0 0 $X=4232000 $Y=560000
X1443 24 1418 mux21_ni $T=4272000 328000 0 0 $X=4272000 $Y=328000
X1444 24 1419 mux21_ni $T=4348000 5664000 1 180 $X=4288000 $Y=5664000
X1445 24 1420 mux21_ni $T=4304000 2184000 0 0 $X=4304000 $Y=2184000
X1446 24 1421 mux21_ni $T=4312000 3344000 0 0 $X=4312000 $Y=3344000
X1447 24 1422 mux21_ni $T=4372000 11232000 1 180 $X=4312000 $Y=11232000
X1448 24 1423 mux21_ni $T=4328000 8912000 0 0 $X=4328000 $Y=8912000
X1449 24 1424 mux21_ni $T=4336000 8448000 0 0 $X=4336000 $Y=8448000
X1450 24 1425 mux21_ni $T=4412000 13088000 1 180 $X=4352000 $Y=13088000
X1451 24 1426 mux21_ni $T=4376000 4040000 0 0 $X=4376000 $Y=4040000
X1452 24 1427 mux21_ni $T=4384000 7288000 0 0 $X=4384000 $Y=7288000
X1453 24 1428 mux21_ni $T=4392000 1024000 0 0 $X=4392000 $Y=1024000
X1454 24 1429 mux21_ni $T=4408000 5664000 0 0 $X=4408000 $Y=5664000
X1455 24 1430 mux21_ni $T=4408000 11696000 0 0 $X=4408000 $Y=11696000
X1456 24 1431 mux21_ni $T=4416000 11000000 0 0 $X=4416000 $Y=11000000
X1457 24 1432 mux21_ni $T=4432000 3576000 0 0 $X=4432000 $Y=3576000
X1458 24 1433 mux21_ni $T=4440000 4040000 0 0 $X=4440000 $Y=4040000
X1459 24 1434 mux21_ni $T=4500000 6128000 1 180 $X=4440000 $Y=6128000
X1460 24 1435 mux21_ni $T=4448000 1720000 0 0 $X=4448000 $Y=1720000
X1461 24 1436 mux21_ni $T=4456000 2416000 0 0 $X=4456000 $Y=2416000
X1462 24 1437 mux21_ni $T=4456000 2648000 0 0 $X=4456000 $Y=2648000
X1463 24 1438 mux21_ni $T=4456000 5200000 0 0 $X=4456000 $Y=5200000
X1464 24 1439 mux21_ni $T=4464000 6824000 0 0 $X=4464000 $Y=6824000
X1465 24 1440 mux21_ni $T=4524000 10536000 1 180 $X=4464000 $Y=10536000
X1466 24 1441 mux21_ni $T=4472000 10768000 0 0 $X=4472000 $Y=10768000
X1467 24 1442 mux21_ni $T=4472000 11928000 0 0 $X=4472000 $Y=11928000
X1468 24 1443 mux21_ni $T=4472000 13088000 0 0 $X=4472000 $Y=13088000
X1469 24 1444 mux21_ni $T=4472000 13320000 0 0 $X=4472000 $Y=13320000
X1470 24 1445 mux21_ni $T=4488000 3112000 0 0 $X=4488000 $Y=3112000
X1471 24 1446 mux21_ni $T=4496000 328000 0 0 $X=4496000 $Y=328000
X1472 24 1447 mux21_ni $T=4496000 1488000 0 0 $X=4496000 $Y=1488000
X1473 24 1448 mux21_ni $T=4496000 9608000 0 0 $X=4496000 $Y=9608000
X1474 24 1449 mux21_ni $T=4520000 96000 0 0 $X=4520000 $Y=96000
X1475 24 1450 mux21_ni $T=4528000 12624000 0 0 $X=4528000 $Y=12624000
X1476 24 1451 mux21_ni $T=4536000 6128000 0 0 $X=4536000 $Y=6128000
X1477 24 1452 mux21_ni $T=4596000 11464000 1 180 $X=4536000 $Y=11464000
X1478 24 1453 mux21_ni $T=4536000 12856000 0 0 $X=4536000 $Y=12856000
X1479 24 1454 mux21_ni $T=4552000 13320000 0 0 $X=4552000 $Y=13320000
X1480 24 1455 mux21_ni $T=4560000 9144000 0 0 $X=4560000 $Y=9144000
X1481 24 1456 mux21_ni $T=4600000 10072000 0 0 $X=4600000 $Y=10072000
X1482 24 1457 mux21_ni $T=4640000 8912000 0 0 $X=4640000 $Y=8912000
X1483 24 1458 mux21_ni $T=4648000 4968000 0 0 $X=4648000 $Y=4968000
X1484 24 1459 mux21_ni $T=4664000 9376000 0 0 $X=4664000 $Y=9376000
X1485 24 1460 mux21_ni $T=4672000 9840000 0 0 $X=4672000 $Y=9840000
X1486 24 1461 mux21_ni $T=4680000 6360000 0 0 $X=4680000 $Y=6360000
X1487 24 1462 mux21_ni $T=4688000 7056000 0 0 $X=4688000 $Y=7056000
X1488 24 1463 mux21_ni $T=4696000 11464000 0 0 $X=4696000 $Y=11464000
X1489 24 1464 mux21_ni $T=4696000 12160000 0 0 $X=4696000 $Y=12160000
X1490 24 1465 mux21_ni $T=4780000 1488000 1 180 $X=4720000 $Y=1488000
X1491 24 1466 mux21_ni $T=4780000 11696000 1 180 $X=4720000 $Y=11696000
X1492 24 1467 mux21_ni $T=4736000 1024000 0 0 $X=4736000 $Y=1024000
X1493 24 1468 mux21_ni $T=4736000 7288000 0 0 $X=4736000 $Y=7288000
X1494 24 1469 mux21_ni $T=4744000 6360000 0 0 $X=4744000 $Y=6360000
X1495 24 1470 mux21_ni $T=4752000 1720000 0 0 $X=4752000 $Y=1720000
X1496 24 1471 mux21_ni $T=4752000 2648000 0 0 $X=4752000 $Y=2648000
X1497 24 1472 mux21_ni $T=4760000 560000 0 0 $X=4760000 $Y=560000
X1498 24 1473 mux21_ni $T=4768000 7520000 0 0 $X=4768000 $Y=7520000
X1499 24 1474 mux21_ni $T=4768000 8680000 0 0 $X=4768000 $Y=8680000
X1500 24 1475 mux21_ni $T=4768000 8912000 0 0 $X=4768000 $Y=8912000
X1501 24 1476 mux21_ni $T=4776000 328000 0 0 $X=4776000 $Y=328000
X1502 24 1477 mux21_ni $T=4784000 4040000 0 0 $X=4784000 $Y=4040000
X1503 24 1478 mux21_ni $T=4808000 1488000 0 0 $X=4808000 $Y=1488000
X1504 24 1479 mux21_ni $T=4816000 2184000 0 0 $X=4816000 $Y=2184000
X1505 24 1480 mux21_ni $T=4816000 5432000 0 0 $X=4816000 $Y=5432000
X1506 24 1481 mux21_ni $T=4816000 12856000 0 0 $X=4816000 $Y=12856000
X1507 24 1482 mux21_ni $T=4824000 6592000 0 0 $X=4824000 $Y=6592000
X1508 24 1483 mux21_ni $T=4856000 13320000 0 0 $X=4856000 $Y=13320000
X1509 24 1484 mux21_ni $T=5052000 5432000 1 180 $X=4992000 $Y=5432000
X1510 24 1485 mux21_ni $T=4992000 7056000 0 0 $X=4992000 $Y=7056000
X1511 24 1486 mux21_ni $T=5000000 13552000 0 0 $X=5000000 $Y=13552000
X1512 24 1487 mux21_ni $T=5016000 4504000 0 0 $X=5016000 $Y=4504000
X1513 24 1488 mux21_ni $T=5076000 12392000 1 180 $X=5016000 $Y=12392000
X1514 24 1489 mux21_ni $T=5076000 12624000 1 180 $X=5016000 $Y=12624000
X1515 24 1490 mux21_ni $T=5100000 11232000 1 180 $X=5040000 $Y=11232000
X1516 24 1491 mux21_ni $T=5108000 8216000 1 180 $X=5048000 $Y=8216000
X1517 24 1492 mux21_ni $T=5072000 7520000 0 0 $X=5072000 $Y=7520000
X1518 24 1493 mux21_ni $T=5080000 9608000 0 0 $X=5080000 $Y=9608000
X1519 24 1494 mux21_ni $T=5096000 1720000 0 0 $X=5096000 $Y=1720000
X1520 24 1495 mux21_ni $T=5128000 6592000 0 0 $X=5128000 $Y=6592000
X1521 24 1496 mux21_ni $T=5152000 4272000 0 0 $X=5152000 $Y=4272000
X1522 24 1497 mux21_ni $T=5160000 3808000 0 0 $X=5160000 $Y=3808000
X1523 24 1498 mux21_ni $T=5176000 1256000 0 0 $X=5176000 $Y=1256000
X1524 24 1499 mux21_ni $T=5236000 3576000 1 180 $X=5176000 $Y=3576000
X1525 24 1500 mux21_ni $T=5192000 8448000 0 0 $X=5192000 $Y=8448000
X1526 24 1501 mux21_ni $T=5200000 328000 0 0 $X=5200000 $Y=328000
X1527 24 1502 mux21_ni $T=5200000 4968000 0 0 $X=5200000 $Y=4968000
X1528 24 1503 mux21_ni $T=5208000 6824000 0 0 $X=5208000 $Y=6824000
X1529 24 1504 mux21_ni $T=5224000 4736000 0 0 $X=5224000 $Y=4736000
X1530 24 1505 mux21_ni $T=5240000 11696000 0 0 $X=5240000 $Y=11696000
X1531 24 1506 mux21_ni $T=5316000 5664000 1 180 $X=5256000 $Y=5664000
X1532 24 1507 mux21_ni $T=5272000 2416000 0 0 $X=5272000 $Y=2416000
X1533 24 1508 mux21_ni $T=5280000 10072000 0 0 $X=5280000 $Y=10072000
X1534 24 1509 mux21_ni $T=5288000 560000 0 0 $X=5288000 $Y=560000
X1535 24 1510 mux21_ni $T=5288000 11464000 0 0 $X=5288000 $Y=11464000
X1536 24 1511 mux21_ni $T=5304000 2880000 0 0 $X=5304000 $Y=2880000
X1537 24 1512 mux21_ni $T=5336000 9840000 0 0 $X=5336000 $Y=9840000
X1538 24 1513 mux21_ni $T=5336000 12160000 0 0 $X=5336000 $Y=12160000
X1539 24 1514 mux21_ni $T=5344000 3112000 0 0 $X=5344000 $Y=3112000
X1540 24 1515 mux21_ni $T=5344000 10536000 0 0 $X=5344000 $Y=10536000
X1541 24 1516 mux21_ni $T=5344000 12392000 0 0 $X=5344000 $Y=12392000
X1542 24 1517 mux21_ni $T=5368000 2648000 0 0 $X=5368000 $Y=2648000
X1543 24 1518 mux21_ni $T=5376000 1720000 0 0 $X=5376000 $Y=1720000
X1544 24 1519 mux21_ni $T=5376000 8680000 0 0 $X=5376000 $Y=8680000
X1545 24 1520 mux21_ni $T=5376000 8912000 0 0 $X=5376000 $Y=8912000
X1546 24 1521 mux21_ni $T=5452000 13320000 1 180 $X=5392000 $Y=13320000
X1547 24 1522 mux21_ni $T=5408000 11000000 0 0 $X=5408000 $Y=11000000
X1548 24 1523 mux21_ni $T=5416000 792000 0 0 $X=5416000 $Y=792000
X1549 24 1524 mux21_ni $T=5416000 8216000 0 0 $X=5416000 $Y=8216000
X1550 24 1525 mux21_ni $T=5424000 1024000 0 0 $X=5424000 $Y=1024000
X1551 24 1526 mux21_ni $T=5424000 12624000 0 0 $X=5424000 $Y=12624000
X1552 24 1527 mux21_ni $T=5448000 96000 0 0 $X=5448000 $Y=96000
X1553 24 1528 mux21_ni $T=5448000 1952000 0 0 $X=5448000 $Y=1952000
X1554 24 1529 mux21_ni $T=5456000 4272000 0 0 $X=5456000 $Y=4272000
X1555 24 1530 mux21_ni $T=5464000 3344000 0 0 $X=5464000 $Y=3344000
X1556 24 1531 mux21_ni $T=5464000 3808000 0 0 $X=5464000 $Y=3808000
X1557 24 1532 mux21_ni $T=5464000 4040000 0 0 $X=5464000 $Y=4040000
X1558 24 1533 mux21_ni $T=5488000 1256000 0 0 $X=5488000 $Y=1256000
X1559 24 1534 mux21_ni $T=5496000 560000 0 0 $X=5496000 $Y=560000
X1560 24 1535 mux21_ni $T=5552000 13320000 0 0 $X=5552000 $Y=13320000
X1561 24 1536 mux21_ni $T=5576000 12856000 0 0 $X=5576000 $Y=12856000
X1562 24 1537 mux21_ni $T=5584000 13088000 0 0 $X=5584000 $Y=13088000
X1563 24 1538 mux21_ni $T=5600000 10304000 0 0 $X=5600000 $Y=10304000
X1564 24 1539 mux21_ni $T=5668000 5432000 1 180 $X=5608000 $Y=5432000
X1565 24 1540 mux21_ni $T=5616000 6128000 0 0 $X=5616000 $Y=6128000
X1566 24 1541 mux21_ni $T=5616000 11928000 0 0 $X=5616000 $Y=11928000
X1567 24 1542 mux21_ni $T=5692000 7056000 1 180 $X=5632000 $Y=7056000
X1568 24 1543 mux21_ni $T=5648000 7984000 0 0 $X=5648000 $Y=7984000
X1569 24 1544 mux21_ni $T=5672000 5432000 0 0 $X=5672000 $Y=5432000
X1570 24 1545 mux21_ni $T=5680000 11928000 0 0 $X=5680000 $Y=11928000
X1571 24 1546 mux21_ni $T=5688000 7752000 0 0 $X=5688000 $Y=7752000
X1572 24 1547 mux21_ni $T=5688000 8680000 0 0 $X=5688000 $Y=8680000
X1573 24 1548 mux21_ni $T=5748000 9840000 1 180 $X=5688000 $Y=9840000
X1574 24 1549 mux21_ni $T=5704000 3808000 0 0 $X=5704000 $Y=3808000
X1575 24 1550 mux21_ni $T=5704000 10536000 0 0 $X=5704000 $Y=10536000
X1576 24 1551 mux21_ni $T=5728000 9376000 0 0 $X=5728000 $Y=9376000
X1577 24 1552 mux21_ni $T=5736000 5432000 0 0 $X=5736000 $Y=5432000
X1578 24 1553 mux21_ni $T=5744000 96000 0 0 $X=5744000 $Y=96000
X1579 24 1554 mux21_ni $T=5744000 12392000 0 0 $X=5744000 $Y=12392000
X1580 24 1555 mux21_ni $T=5760000 1952000 0 0 $X=5760000 $Y=1952000
X1581 24 1556 mux21_ni $T=5760000 2184000 0 0 $X=5760000 $Y=2184000
X1582 24 1557 mux21_ni $T=5760000 4504000 0 0 $X=5760000 $Y=4504000
X1583 24 1558 mux21_ni $T=5820000 6360000 1 180 $X=5760000 $Y=6360000
X1584 24 1559 mux21_ni $T=5760000 13552000 0 0 $X=5760000 $Y=13552000
X1585 24 1560 mux21_ni $T=5800000 560000 0 0 $X=5800000 $Y=560000
X1586 24 1561 mux21_ni $T=5800000 9144000 0 0 $X=5800000 $Y=9144000
X1587 24 1562 mux21_ni $T=5816000 6824000 0 0 $X=5816000 $Y=6824000
X1588 24 1563 mux21_ni $T=5824000 6360000 0 0 $X=5824000 $Y=6360000
X1589 24 1564 mux21_ni $T=5840000 9840000 0 0 $X=5840000 $Y=9840000
X1590 24 1565 mux21_ni $T=5872000 328000 0 0 $X=5872000 $Y=328000
X1591 24 1566 mux21_ni $T=5872000 8448000 0 0 $X=5872000 $Y=8448000
X1592 24 1567 mux21_ni $T=5904000 13088000 0 0 $X=5904000 $Y=13088000
X1593 24 1568 mux21_ni $T=5936000 3112000 0 0 $X=5936000 $Y=3112000
X1594 24 1569 mux21_ni $T=6004000 7288000 1 180 $X=5944000 $Y=7288000
X1595 24 1570 mux21_ni $T=5968000 4736000 0 0 $X=5968000 $Y=4736000
X1596 24 1571 mux21_ni $T=5968000 7056000 0 0 $X=5968000 $Y=7056000
X1597 24 1572 mux21_ni $T=5976000 3576000 0 0 $X=5976000 $Y=3576000
X1598 24 1573 mux21_ni $T=5984000 2648000 0 0 $X=5984000 $Y=2648000
X1599 24 1574 mux21_ni $T=5984000 4272000 0 0 $X=5984000 $Y=4272000
X1600 24 1575 mux21_ni $T=5992000 8912000 0 0 $X=5992000 $Y=8912000
X1601 24 1576 mux21_ni $T=6000000 8216000 0 0 $X=6000000 $Y=8216000
X1602 24 1577 mux21_ni $T=6000000 11464000 0 0 $X=6000000 $Y=11464000
X1603 24 1578 mux21_ni $T=6016000 3344000 0 0 $X=6016000 $Y=3344000
X1604 24 1579 mux21_ni $T=6024000 7984000 0 0 $X=6024000 $Y=7984000
X1605 24 1580 mux21_ni $T=6032000 2880000 0 0 $X=6032000 $Y=2880000
X1606 24 1581 mux21_ni $T=6040000 1256000 0 0 $X=6040000 $Y=1256000
X1607 24 1582 mux21_ni $T=6048000 2416000 0 0 $X=6048000 $Y=2416000
X1608 24 1583 mux21_ni $T=6056000 8912000 0 0 $X=6056000 $Y=8912000
X1609 24 1584 mux21_ni $T=6056000 11000000 0 0 $X=6056000 $Y=11000000
X1610 24 1585 mux21_ni $T=6064000 1024000 0 0 $X=6064000 $Y=1024000
X1611 24 1586 mux21_ni $T=6064000 7288000 0 0 $X=6064000 $Y=7288000
X1612 24 1587 mux21_ni $T=6072000 2184000 0 0 $X=6072000 $Y=2184000
X1613 24 1588 mux21_ni $T=6080000 792000 0 0 $X=6080000 $Y=792000
X1614 24 1589 mux21_ni $T=6080000 11232000 0 0 $X=6080000 $Y=11232000
X1615 24 1590 mux21_ni $T=6080000 11696000 0 0 $X=6080000 $Y=11696000
X1616 24 1591 mux21_ni $T=6088000 11928000 0 0 $X=6088000 $Y=11928000
X1617 24 1592 mux21_ni $T=6088000 12160000 0 0 $X=6088000 $Y=12160000
X1618 24 1593 mux21_ni $T=6104000 560000 0 0 $X=6104000 $Y=560000
X1619 24 1594 mux21_ni $T=6120000 8912000 0 0 $X=6120000 $Y=8912000
X1620 24 1595 mux21_ni $T=6128000 10768000 0 0 $X=6128000 $Y=10768000
X1621 24 1596 mux21_ni $T=6128000 12392000 0 0 $X=6128000 $Y=12392000
X1622 24 1597 mux21_ni $T=6128000 12624000 0 0 $X=6128000 $Y=12624000
X1623 24 1598 mux21_ni $T=6144000 9840000 0 0 $X=6144000 $Y=9840000
X1624 24 1599 mux21_ni $T=6160000 10536000 0 0 $X=6160000 $Y=10536000
X1625 24 1600 mux21_ni $T=6184000 10304000 0 0 $X=6184000 $Y=10304000
X1626 24 1601 mux21_ni $T=6256000 3808000 0 0 $X=6256000 $Y=3808000
X1627 24 1602 mux21_ni $T=6256000 13552000 0 0 $X=6256000 $Y=13552000
X1628 24 1603 mux21_ni $T=6264000 4040000 0 0 $X=6264000 $Y=4040000
X1629 24 1604 mux21_ni $T=6324000 5432000 1 180 $X=6264000 $Y=5432000
X1630 24 1605 mux21_ni $T=6280000 3576000 0 0 $X=6280000 $Y=3576000
X1631 24 1606 mux21_ni $T=6280000 4736000 0 0 $X=6280000 $Y=4736000
X1632 24 1607 mux21_ni $T=6296000 4272000 0 0 $X=6296000 $Y=4272000
X1633 24 1608 mux21_ni $T=6296000 11464000 0 0 $X=6296000 $Y=11464000
X1634 24 1609 mux21_ni $T=6328000 5432000 0 0 $X=6328000 $Y=5432000
X1635 24 1610 mux21_ni $T=6328000 12856000 0 0 $X=6328000 $Y=12856000
X1636 24 1611 mux21_ni $T=6336000 8448000 0 0 $X=6336000 $Y=8448000
X1637 24 1612 mux21_ni $T=6336000 11696000 0 0 $X=6336000 $Y=11696000
X1638 24 1613 mux21_ni $T=6344000 11000000 0 0 $X=6344000 $Y=11000000
X1639 24 1614 mux21_ni $T=6352000 13320000 0 0 $X=6352000 $Y=13320000
X1640 24 1615 mux21_ni $T=6360000 1488000 0 0 $X=6360000 $Y=1488000
X1641 24 1616 mux21_ni $T=6360000 4272000 0 0 $X=6360000 $Y=4272000
X1642 24 1617 mux21_ni $T=6368000 7984000 0 0 $X=6368000 $Y=7984000
X1643 24 1618 mux21_ni $T=6368000 11928000 0 0 $X=6368000 $Y=11928000
X1644 24 1619 mux21_ni $T=6376000 1024000 0 0 $X=6376000 $Y=1024000
X1645 24 1620 mux21_ni $T=6392000 9608000 0 0 $X=6392000 $Y=9608000
X1646 24 1621 mux21_ni $T=6460000 6824000 1 180 $X=6400000 $Y=6824000
X1647 24 1622 mux21_ni $T=6416000 792000 0 0 $X=6416000 $Y=792000
X1648 24 1623 mux21_ni $T=6416000 2416000 0 0 $X=6416000 $Y=2416000
X1649 24 1624 mux21_ni $T=6432000 1720000 0 0 $X=6432000 $Y=1720000
X1650 24 1625 mux21_ni $T=6440000 1952000 0 0 $X=6440000 $Y=1952000
X1651 24 1626 mux21_ni $T=6440000 3344000 0 0 $X=6440000 $Y=3344000
X1652 24 1627 mux21_ni $T=6440000 12624000 0 0 $X=6440000 $Y=12624000
X1653 24 1628 mux21_ni $T=6440000 13088000 0 0 $X=6440000 $Y=13088000
X1654 24 1629 mux21_ni $T=6516000 7752000 1 180 $X=6456000 $Y=7752000
X1655 24 1630 mux21_ni $T=6472000 10304000 0 0 $X=6472000 $Y=10304000
X1656 24 1631 mux21_ni $T=6520000 7752000 0 0 $X=6520000 $Y=7752000
X1657 24 1632 mux21_ni $T=6588000 6824000 1 180 $X=6528000 $Y=6824000
X1658 24 1633 mux21_ni $T=6528000 8912000 0 0 $X=6528000 $Y=8912000
X1659 24 1634 mux21_ni $T=6536000 8216000 0 0 $X=6536000 $Y=8216000
X1660 24 1635 mux21_ni $T=6552000 328000 0 0 $X=6552000 $Y=328000
X1661 24 1636 mux21_ni $T=6576000 5200000 0 0 $X=6576000 $Y=5200000
X1662 24 1637 mux21_ni $T=6592000 11232000 0 0 $X=6592000 $Y=11232000
X1663 24 1638 mux21_ni $T=6600000 8216000 0 0 $X=6600000 $Y=8216000
X1664 24 1639 mux21_ni $T=6692000 6360000 1 180 $X=6632000 $Y=6360000
X1665 24 1640 mux21_ni $T=6632000 9840000 0 0 $X=6632000 $Y=9840000
X1666 24 1641 mux21_ni $T=6640000 4736000 0 0 $X=6640000 $Y=4736000
X1667 24 1642 mux21_ni $T=6708000 2880000 1 180 $X=6648000 $Y=2880000
X1668 24 1643 mux21_ni $T=6708000 5896000 1 180 $X=6648000 $Y=5896000
X1669 24 1644 mux21_ni $T=6656000 96000 0 0 $X=6656000 $Y=96000
X1670 24 1645 mux21_ni $T=6664000 560000 0 0 $X=6664000 $Y=560000
X1671 24 1646 mux21_ni $T=6672000 4504000 0 0 $X=6672000 $Y=4504000
X1672 24 1647 mux21_ni $T=6680000 8680000 0 0 $X=6680000 $Y=8680000
X1673 24 1648 mux21_ni $T=6688000 10768000 0 0 $X=6688000 $Y=10768000
X1674 24 1649 mux21_ni $T=6736000 4968000 0 0 $X=6736000 $Y=4968000
X1675 24 1650 mux21_ni $T=6736000 10072000 0 0 $X=6736000 $Y=10072000
X1676 24 1651 mux21_ni $T=6744000 3344000 0 0 $X=6744000 $Y=3344000
X1677 24 1652 mux21_ni $T=6768000 1720000 0 0 $X=6768000 $Y=1720000
X1678 24 1653 mux21_ni $T=6776000 1952000 0 0 $X=6776000 $Y=1952000
X1679 24 1654 mux21_ni $T=6784000 8448000 0 0 $X=6784000 $Y=8448000
X1680 24 1655 mux21_ni $T=6800000 2416000 0 0 $X=6800000 $Y=2416000
X1681 24 1656 mux21_ni $T=6800000 3576000 0 0 $X=6800000 $Y=3576000
X1682 24 1657 mux21_ni $T=6824000 2880000 0 0 $X=6824000 $Y=2880000
X1683 24 1658 mux21_ni $T=6832000 5664000 0 0 $X=6832000 $Y=5664000
X1684 24 1659 mux21_ni $T=6848000 7056000 0 0 $X=6848000 $Y=7056000
X1685 24 1660 mux21_ni $T=6880000 12856000 0 0 $X=6880000 $Y=12856000
X1686 24 1661 mux21_ni $T=6940000 13320000 1 180 $X=6880000 $Y=13320000
X1687 24 1662 mux21_ni $T=6948000 12160000 1 180 $X=6888000 $Y=12160000
X1688 24 1663 mux21_ni $T=6896000 6824000 0 0 $X=6896000 $Y=6824000
X1689 24 1664 mux21_ni $T=6896000 8216000 0 0 $X=6896000 $Y=8216000
X1690 24 1665 mux21_ni $T=6912000 13088000 0 0 $X=6912000 $Y=13088000
X1691 24 1666 mux21_ni $T=6920000 4736000 0 0 $X=6920000 $Y=4736000
X1692 24 1667 mux21_ni $T=6928000 2184000 0 0 $X=6928000 $Y=2184000
X1693 24 1668 mux21_ni $T=6936000 7984000 0 0 $X=6936000 $Y=7984000
X1694 24 1669 mux21_ni $T=6944000 5432000 0 0 $X=6944000 $Y=5432000
X1695 24 1670 mux21_ni $T=6960000 5896000 0 0 $X=6960000 $Y=5896000
X1696 24 1671 mux21_ni $T=6960000 8680000 0 0 $X=6960000 $Y=8680000
X1697 24 1672 mux21_ni $T=6976000 13320000 0 0 $X=6976000 $Y=13320000
X1698 24 1673 mux21_ni $T=6984000 1024000 0 0 $X=6984000 $Y=1024000
X1699 24 1674 mux21_ni $T=6992000 10768000 0 0 $X=6992000 $Y=10768000
X1700 24 1675 mux21_ni $T=7000000 6128000 0 0 $X=7000000 $Y=6128000
X1701 24 1676 mux21_ni $T=7000000 7984000 0 0 $X=7000000 $Y=7984000
X1702 24 1677 mux21_ni $T=7016000 11000000 0 0 $X=7016000 $Y=11000000
X1703 24 1678 mux21_ni $T=7024000 3344000 0 0 $X=7024000 $Y=3344000
X1704 24 1679 mux21_ni $T=7024000 8680000 0 0 $X=7024000 $Y=8680000
X1705 24 1680 mux21_ni $T=7048000 12392000 0 0 $X=7048000 $Y=12392000
X1706 24 1681 mux21_ni $T=7072000 4040000 0 0 $X=7072000 $Y=4040000
X1707 24 1682 mux21_ni $T=7080000 2648000 0 0 $X=7080000 $Y=2648000
X1708 24 1683 mux21_ni $T=7172000 3112000 1 180 $X=7112000 $Y=3112000
X1709 24 1684 mux21_ni $T=7136000 10536000 0 0 $X=7136000 $Y=10536000
X1710 24 1685 mux21_ni $T=7160000 3576000 0 0 $X=7160000 $Y=3576000
X1711 24 1686 mux21_ni $T=7244000 6592000 1 180 $X=7184000 $Y=6592000
X1712 24 1687 mux21_ni $T=7192000 1488000 0 0 $X=7192000 $Y=1488000
X1713 24 1688 mux21_ni $T=7252000 9376000 1 180 $X=7192000 $Y=9376000
X1714 24 1689 mux21_ni $T=7200000 10304000 0 0 $X=7200000 $Y=10304000
X1715 24 1690 mux21_ni $T=7208000 3112000 0 0 $X=7208000 $Y=3112000
X1716 24 1691 mux21_ni $T=7224000 6360000 0 0 $X=7224000 $Y=6360000
X1717 24 1692 mux21_ni $T=7240000 12624000 0 0 $X=7240000 $Y=12624000
X1718 24 1693 mux21_ni $T=7300000 12856000 1 180 $X=7240000 $Y=12856000
X1719 24 1694 mux21_ni $T=7248000 6592000 0 0 $X=7248000 $Y=6592000
X1720 24 1695 mux21_ni $T=7316000 10072000 1 180 $X=7256000 $Y=10072000
X1721 24 1696 mux21_ni $T=7280000 560000 0 0 $X=7280000 $Y=560000
X1722 24 1697 mux21_ni $T=7340000 4736000 1 180 $X=7280000 $Y=4736000
X1723 24 1698 mux21_ni $T=7288000 6360000 0 0 $X=7288000 $Y=6360000
X1724 24 1699 mux21_ni $T=7328000 1256000 0 0 $X=7328000 $Y=1256000
X1725 24 1700 mux21_ni $T=7388000 7056000 1 180 $X=7328000 $Y=7056000
X1726 24 1701 mux21_ni $T=7336000 8448000 0 0 $X=7336000 $Y=8448000
X1727 24 1702 mux21_ni $T=7344000 11464000 0 0 $X=7344000 $Y=11464000
X1728 24 1703 mux21_ni $T=7344000 11696000 0 0 $X=7344000 $Y=11696000
X1729 24 1704 mux21_ni $T=7352000 10768000 0 0 $X=7352000 $Y=10768000
X1730 24 1705 mux21_ni $T=7384000 3344000 0 0 $X=7384000 $Y=3344000
X1731 24 1706 mux21_ni $T=7476000 8216000 1 180 $X=7416000 $Y=8216000
X1732 24 1707 mux21_ni $T=7492000 9608000 1 180 $X=7432000 $Y=9608000
X1733 24 1708 mux21_ni $T=7508000 7752000 1 180 $X=7448000 $Y=7752000
X1734 24 1709 mux21_ni $T=7448000 11232000 0 0 $X=7448000 $Y=11232000
X1735 24 1710 mux21_ni $T=7464000 7288000 0 0 $X=7464000 $Y=7288000
X1736 24 1711 mux21_ni $T=7472000 5432000 0 0 $X=7472000 $Y=5432000
X1737 24 1712 mux21_ni $T=7480000 3344000 0 0 $X=7480000 $Y=3344000
X1738 24 1713 mux21_ni $T=7556000 328000 1 180 $X=7496000 $Y=328000
X1739 24 1714 mux21_ni $T=7512000 3112000 0 0 $X=7512000 $Y=3112000
X1740 24 1715 mux21_ni $T=7512000 7752000 0 0 $X=7512000 $Y=7752000
X1741 24 1716 mux21_ni $T=7520000 792000 0 0 $X=7520000 $Y=792000
X1742 24 1717 mux21_ni $T=7528000 9608000 0 0 $X=7528000 $Y=9608000
X1743 24 1718 mux21_ni $T=7536000 4272000 0 0 $X=7536000 $Y=4272000
X1744 24 1719 mux21_ni $T=7536000 8216000 0 0 $X=7536000 $Y=8216000
X1745 24 1720 mux21_ni $T=7612000 11000000 1 180 $X=7552000 $Y=11000000
X1746 24 1721 mux21_ni $T=7568000 10072000 0 0 $X=7568000 $Y=10072000
X1747 24 1722 mux21_ni $T=7592000 4736000 0 0 $X=7592000 $Y=4736000
X1748 24 1723 mux21_ni $T=7592000 9840000 0 0 $X=7592000 $Y=9840000
X1749 24 1724 mux21_ni $T=7600000 4272000 0 0 $X=7600000 $Y=4272000
X1750 24 1725 mux21_ni $T=7600000 8216000 0 0 $X=7600000 $Y=8216000
X1751 24 1726 mux21_ni $T=7600000 9144000 0 0 $X=7600000 $Y=9144000
X1752 24 1727 mux21_ni $T=7600000 9376000 0 0 $X=7600000 $Y=9376000
X1753 24 1728 mux21_ni $T=7616000 328000 0 0 $X=7616000 $Y=328000
X1754 24 1729 mux21_ni $T=7616000 11000000 0 0 $X=7616000 $Y=11000000
X1755 24 1730 mux21_ni $T=7692000 1952000 1 180 $X=7632000 $Y=1952000
X1756 24 1731 mux21_ni $T=7640000 2416000 0 0 $X=7640000 $Y=2416000
X1757 24 1732 mux21_ni $T=7648000 13320000 0 0 $X=7648000 $Y=13320000
X1758 24 1733 mux21_ni $T=7664000 3808000 0 0 $X=7664000 $Y=3808000
X1759 24 1734 mux21_ni $T=7724000 10768000 1 180 $X=7664000 $Y=10768000
X1760 24 1735 mux21_ni $T=7680000 96000 0 0 $X=7680000 $Y=96000
X1761 24 1736 mux21_ni $T=7680000 8680000 0 0 $X=7680000 $Y=8680000
X1762 24 1737 mux21_ni $T=7696000 1952000 0 0 $X=7696000 $Y=1952000
X1763 24 1738 mux21_ni $T=7704000 6128000 0 0 $X=7704000 $Y=6128000
X1764 24 1739 mux21_ni $T=7704000 8912000 0 0 $X=7704000 $Y=8912000
X1765 24 1740 mux21_ni $T=7712000 3576000 0 0 $X=7712000 $Y=3576000
X1766 24 1741 mux21_ni $T=7736000 12856000 0 0 $X=7736000 $Y=12856000
X1767 24 1742 mux21_ni $T=7736000 13320000 0 0 $X=7736000 $Y=13320000
X1768 24 1743 mux21_ni $T=7744000 4040000 0 0 $X=7744000 $Y=4040000
X1769 24 1744 mux21_ni $T=7744000 5896000 0 0 $X=7744000 $Y=5896000
X1770 24 1745 mux21_ni $T=7844000 12160000 1 180 $X=7784000 $Y=12160000
X1771 24 1746 mux21_ni $T=7892000 11464000 1 180 $X=7832000 $Y=11464000
X1772 24 1747 mux21_ni $T=7872000 5200000 0 0 $X=7872000 $Y=5200000
X1773 24 1748 mux21_ni $T=7880000 1256000 0 0 $X=7880000 $Y=1256000
X1774 24 1749 mux21_ni $T=7880000 5432000 0 0 $X=7880000 $Y=5432000
X1775 24 1750 mux21_ni $T=7940000 8448000 1 180 $X=7880000 $Y=8448000
X1776 24 1751 mux21_ni $T=7936000 11464000 0 0 $X=7936000 $Y=11464000
X1777 24 1752 mux21_ni $T=7944000 8448000 0 0 $X=7944000 $Y=8448000
X1778 24 1753 mux21_ni $T=7952000 560000 0 0 $X=7952000 $Y=560000
X1779 24 1754 mux21_ni $T=8020000 7288000 1 180 $X=7960000 $Y=7288000
X1780 24 1755 mux21_ni $T=8020000 11696000 1 180 $X=7960000 $Y=11696000
X1781 24 1756 mux21_ni $T=8028000 10768000 1 180 $X=7968000 $Y=10768000
X1782 24 1757 mux21_ni $T=7984000 6128000 0 0 $X=7984000 $Y=6128000
X1783 24 1758 mux21_ni $T=7984000 11232000 0 0 $X=7984000 $Y=11232000
X1784 24 1759 mux21_ni $T=8052000 3576000 1 180 $X=7992000 $Y=3576000
X1785 24 1760 mux21_ni $T=8024000 11696000 0 0 $X=8024000 $Y=11696000
X1786 24 1761 mux21_ni $T=8032000 4968000 0 0 $X=8032000 $Y=4968000
X1787 24 1762 mux21_ni $T=8032000 10768000 0 0 $X=8032000 $Y=10768000
X1788 24 1763 mux21_ni $T=8064000 1488000 0 0 $X=8064000 $Y=1488000
X1789 24 1764 mux21_ni $T=8064000 6360000 0 0 $X=8064000 $Y=6360000
X1790 24 1765 mux21_ni $T=8064000 7984000 0 0 $X=8064000 $Y=7984000
X1791 24 1766 mux21_ni $T=8096000 9376000 0 0 $X=8096000 $Y=9376000
X1792 24 1767 mux21_ni $T=8156000 13088000 1 180 $X=8096000 $Y=13088000
X1793 24 1768 mux21_ni $T=8180000 2648000 1 180 $X=8120000 $Y=2648000
X1794 24 1769 mux21_ni $T=8120000 4736000 0 0 $X=8120000 $Y=4736000
X1795 24 1770 mux21_ni $T=8120000 10536000 0 0 $X=8120000 $Y=10536000
X1796 24 1771 mux21_ni $T=8128000 7520000 0 0 $X=8128000 $Y=7520000
X1797 24 1772 mux21_ni $T=8160000 3112000 0 0 $X=8160000 $Y=3112000
X1798 24 1773 mux21_ni $T=8160000 4272000 0 0 $X=8160000 $Y=4272000
X1799 24 1774 mux21_ni $T=8176000 6824000 0 0 $X=8176000 $Y=6824000
X1800 24 1775 mux21_ni $T=8236000 12160000 1 180 $X=8176000 $Y=12160000
X1801 24 1776 mux21_ni $T=8192000 1256000 0 0 $X=8192000 $Y=1256000
X1802 24 1777 mux21_ni $T=8240000 11464000 0 0 $X=8240000 $Y=11464000
X1803 24 1778 mux21_ni $T=8256000 8448000 0 0 $X=8256000 $Y=8448000
X1804 24 1779 mux21_ni $T=8256000 11696000 0 0 $X=8256000 $Y=11696000
X1805 24 1780 mux21_ni $T=8264000 5200000 0 0 $X=8264000 $Y=5200000
X1806 24 1781 mux21_ni $T=8288000 11232000 0 0 $X=8288000 $Y=11232000
X1807 24 1782 mux21_ni $T=8356000 3576000 1 180 $X=8296000 $Y=3576000
X1808 24 1783 mux21_ni $T=8296000 6592000 0 0 $X=8296000 $Y=6592000
X1809 24 1784 mux21_ni $T=8312000 560000 0 0 $X=8312000 $Y=560000
X1810 24 1785 mux21_ni $T=8320000 5664000 0 0 $X=8320000 $Y=5664000
X1811 24 1786 mux21_ni $T=8420000 3808000 1 180 $X=8360000 $Y=3808000
X1812 24 1787 mux21_ni $T=8368000 1488000 0 0 $X=8368000 $Y=1488000
X1813 24 1788 mux21_ni $T=8376000 6128000 0 0 $X=8376000 $Y=6128000
X1814 24 1789 mux21_ni $T=8444000 1952000 1 180 $X=8384000 $Y=1952000
X1815 24 1790 mux21_ni $T=8384000 8680000 0 0 $X=8384000 $Y=8680000
X1816 24 1791 mux21_ni $T=8384000 8912000 0 0 $X=8384000 $Y=8912000
X1817 24 1792 mux21_ni $T=8392000 2416000 0 0 $X=8392000 $Y=2416000
X1818 24 1793 mux21_ni $T=8408000 8216000 0 0 $X=8408000 $Y=8216000
X1819 24 1794 mux21_ni $T=8476000 4968000 1 180 $X=8416000 $Y=4968000
X1820 24 1795 mux21_ni $T=8432000 7520000 0 0 $X=8432000 $Y=7520000
X1821 24 1796 mux21_ni $T=8432000 10304000 0 0 $X=8432000 $Y=10304000
X1822 24 1797 mux21_ni $T=8464000 7752000 0 0 $X=8464000 $Y=7752000
X1823 24 1798 mux21_ni $T=8488000 10536000 0 0 $X=8488000 $Y=10536000
X1824 24 1799 mux21_ni $T=8496000 792000 0 0 $X=8496000 $Y=792000
X1825 24 1800 mux21_ni $T=8496000 1256000 0 0 $X=8496000 $Y=1256000
X1826 24 1801 mux21_ni $T=8496000 4272000 0 0 $X=8496000 $Y=4272000
X1827 24 1802 mux21_ni $T=8512000 6824000 0 0 $X=8512000 $Y=6824000
X1828 24 1803 mux21_ni $T=8544000 5200000 0 0 $X=8544000 $Y=5200000
X1829 24 1804 mux21_ni $T=8560000 5432000 0 0 $X=8560000 $Y=5432000
X1830 24 1805 mux21_ni $T=8568000 4504000 0 0 $X=8568000 $Y=4504000
X1831 24 1806 mux21_ni $T=8568000 11232000 0 0 $X=8568000 $Y=11232000
X1832 24 1807 mux21_ni $T=8584000 5896000 0 0 $X=8584000 $Y=5896000
X1833 24 1808 mux21_ni $T=8592000 3344000 0 0 $X=8592000 $Y=3344000
X1834 24 1809 mux21_ni $T=8592000 4968000 0 0 $X=8592000 $Y=4968000
X1835 24 1810 mux21_ni $T=8600000 6360000 0 0 $X=8600000 $Y=6360000
X1836 24 1811 mux21_ni $T=8660000 11000000 1 180 $X=8600000 $Y=11000000
X1837 24 1812 mux21_ni $T=8624000 10072000 0 0 $X=8624000 $Y=10072000
X1838 24 1813 mux21_ni $T=8648000 5896000 0 0 $X=8648000 $Y=5896000
X1839 24 1814 mux21_ni $T=8672000 1488000 0 0 $X=8672000 $Y=1488000
X1840 24 1815 mux21_ni $T=8680000 2648000 0 0 $X=8680000 $Y=2648000
X1841 24 1816 mux21_ni $T=8680000 4040000 0 0 $X=8680000 $Y=4040000
X1842 24 1817 mux21_ni $T=8688000 328000 0 0 $X=8688000 $Y=328000
X1843 24 1818 mux21_ni $T=8696000 9840000 0 0 $X=8696000 $Y=9840000
X1844 24 1819 mux21_ni $T=8704000 96000 0 0 $X=8704000 $Y=96000
X1845 24 1820 mux21_ni $T=8712000 4968000 0 0 $X=8712000 $Y=4968000
X1846 24 1821 mux21_ni $T=8812000 8448000 1 180 $X=8752000 $Y=8448000
X1847 24 1822 mux21_ni $T=8752000 11000000 0 0 $X=8752000 $Y=11000000
X1848 24 1823 mux21_ni $T=8820000 1952000 1 180 $X=8760000 $Y=1952000
X1849 24 1824 mux21_ni $T=8760000 9840000 0 0 $X=8760000 $Y=9840000
X1850 24 1825 mux21_ni $T=8784000 328000 0 0 $X=8784000 $Y=328000
X1851 24 1826 mux21_ni $T=8792000 10304000 0 0 $X=8792000 $Y=10304000
X1852 24 1827 mux21_ni $T=8792000 10536000 0 0 $X=8792000 $Y=10536000
X1853 24 1828 mux21_ni $T=8800000 792000 0 0 $X=8800000 $Y=792000
X1854 24 1829 mux21_ni $T=8808000 7752000 0 0 $X=8808000 $Y=7752000
X1855 24 1830 mux21_ni $T=8816000 9376000 0 0 $X=8816000 $Y=9376000
X1856 24 1831 mux21_ni $T=8916000 7288000 1 180 $X=8856000 $Y=7288000
X1857 24 1832 mux21_ni $T=8896000 4736000 0 0 $X=8896000 $Y=4736000
X1858 24 1833 mux21_ni $T=8964000 12856000 1 180 $X=8904000 $Y=12856000
X1859 24 1834 mux21_ni $T=8996000 6128000 1 180 $X=8936000 $Y=6128000
X1860 24 1835 mux21_ni $T=8952000 1488000 0 0 $X=8952000 $Y=1488000
X1861 24 1836 mux21_ni $T=8960000 5896000 0 0 $X=8960000 $Y=5896000
X1862 24 1837 mux21_ni $T=8968000 2184000 0 0 $X=8968000 $Y=2184000
X1863 24 1838 mux21_ni $T=8992000 3112000 0 0 $X=8992000 $Y=3112000
X1864 24 1839 mux21_ni $T=8992000 4040000 0 0 $X=8992000 $Y=4040000
X1865 24 1840 mux21_ni $T=9000000 6128000 0 0 $X=9000000 $Y=6128000
X1866 24 1841 mux21_ni $T=9008000 3344000 0 0 $X=9008000 $Y=3344000
X1867 24 1842 mux21_ni $T=9016000 560000 0 0 $X=9016000 $Y=560000
X1868 24 1843 mux21_ni $T=9016000 1720000 0 0 $X=9016000 $Y=1720000
X1869 24 1844 mux21_ni $T=9016000 2880000 0 0 $X=9016000 $Y=2880000
X1870 24 1845 mux21_ni $T=9032000 2184000 0 0 $X=9032000 $Y=2184000
X1871 24 1846 mux21_ni $T=9092000 11232000 1 180 $X=9032000 $Y=11232000
X1872 24 1847 mux21_ni $T=9048000 1256000 0 0 $X=9048000 $Y=1256000
X1873 24 1848 mux21_ni $T=9116000 1024000 1 180 $X=9056000 $Y=1024000
X1874 24 1849 mux21_ni $T=9056000 9144000 0 0 $X=9056000 $Y=9144000
X1875 24 1850 mux21_ni $T=9056000 11696000 0 0 $X=9056000 $Y=11696000
X1876 24 1851 mux21_ni $T=9132000 11464000 1 180 $X=9072000 $Y=11464000
X1877 24 1852 mux21_ni $T=9096000 2184000 0 0 $X=9096000 $Y=2184000
X1878 24 1853 mux21_ni $T=9096000 3576000 0 0 $X=9096000 $Y=3576000
X1879 24 1854 mux21_ni $T=9104000 1952000 0 0 $X=9104000 $Y=1952000
X1880 24 1855 mux21_ni $T=9112000 8216000 0 0 $X=9112000 $Y=8216000
X1881 24 1856 mux21_ni $T=9120000 8448000 0 0 $X=9120000 $Y=8448000
X1882 24 1857 mux21_ni $T=9120000 9376000 0 0 $X=9120000 $Y=9376000
X1883 24 1858 mux21_ni $T=9136000 5432000 0 0 $X=9136000 $Y=5432000
X1884 24 1859 mux21_ni $T=9144000 328000 0 0 $X=9144000 $Y=328000
X1885 24 1860 mux21_ni $T=9160000 3576000 0 0 $X=9160000 $Y=3576000
X1886 24 1861 mux21_ni $T=9160000 4272000 0 0 $X=9160000 $Y=4272000
X1887 24 1862 mux21_ni $T=9168000 7056000 0 0 $X=9168000 $Y=7056000
X1888 24 1863 mux21_ni $T=9168000 11928000 0 0 $X=9168000 $Y=11928000
X1889 24 1864 mux21_ni $T=9236000 7984000 1 180 $X=9176000 $Y=7984000
X1890 24 1865 mux21_ni $T=9236000 12160000 1 180 $X=9176000 $Y=12160000
X1891 24 1866 mux21_ni $T=9184000 10304000 0 0 $X=9184000 $Y=10304000
X1892 24 1867 mux21_ni $T=9192000 10768000 0 0 $X=9192000 $Y=10768000
X1893 24 1868 mux21_ni $T=9260000 13320000 1 180 $X=9200000 $Y=13320000
X1894 24 1869 mux21_ni $T=9208000 9840000 0 0 $X=9208000 $Y=9840000
X1895 24 1870 mux21_ni $T=9208000 10536000 0 0 $X=9208000 $Y=10536000
X1896 24 1871 mux21_ni $T=9232000 1488000 0 0 $X=9232000 $Y=1488000
X1897 24 1872 mux21_ni $T=9292000 5664000 1 180 $X=9232000 $Y=5664000
X1898 24 1873 mux21_ni $T=9232000 8912000 0 0 $X=9232000 $Y=8912000
X1899 24 1874 mux21_ni $T=9232000 11232000 0 0 $X=9232000 $Y=11232000
X1900 24 1875 mux21_ni $T=9256000 6360000 0 0 $X=9256000 $Y=6360000
X1901 24 1876 mux21_ni $T=9256000 10768000 0 0 $X=9256000 $Y=10768000
X1902 24 1877 mux21_ni $T=9264000 4736000 0 0 $X=9264000 $Y=4736000
X1903 24 1878 mux21_ni $T=9264000 5896000 0 0 $X=9264000 $Y=5896000
X1904 24 1879 mux21_ni $T=9356000 3112000 1 180 $X=9296000 $Y=3112000
X1905 24 1880 mux21_ni $T=9356000 7984000 1 180 $X=9296000 $Y=7984000
X1906 24 1881 mux21_ni $T=9304000 6128000 0 0 $X=9304000 $Y=6128000
X1907 24 1882 mux21_ni $T=9312000 3344000 0 0 $X=9312000 $Y=3344000
X1908 24 1883 mux21_ni $T=9320000 1720000 0 0 $X=9320000 $Y=1720000
X1909 24 1884 mux21_ni $T=9328000 9840000 0 0 $X=9328000 $Y=9840000
X1910 24 1885 mux21_ni $T=9344000 5200000 0 0 $X=9344000 $Y=5200000
X1911 24 1886 mux21_ni $T=9352000 5664000 0 0 $X=9352000 $Y=5664000
X1912 24 1887 mux21_ni $T=9360000 3112000 0 0 $X=9360000 $Y=3112000
X1913 24 1888 mux21_ni $T=9376000 3344000 0 0 $X=9376000 $Y=3344000
X1914 24 1889 mux21_ni $T=9460000 2184000 1 180 $X=9400000 $Y=2184000
X1915 24 1890 mux21_ni $T=9416000 1256000 0 0 $X=9416000 $Y=1256000
X1916 24 1891 mux21_ni $T=9448000 328000 0 0 $X=9448000 $Y=328000
X1917 24 1892 mux21_ni $T=9456000 2648000 0 0 $X=9456000 $Y=2648000
X1918 24 1893 mux21_ni $T=9472000 7056000 0 0 $X=9472000 $Y=7056000
X1919 24 1894 mux21_ni $T=9480000 4968000 0 0 $X=9480000 $Y=4968000
X1920 24 1895 mux21_ni $T=9496000 2184000 0 0 $X=9496000 $Y=2184000
X1921 24 1896 mux21_ni $T=9504000 96000 0 0 $X=9504000 $Y=96000
X1922 24 1897 mux21_ni $T=9560000 3808000 0 0 $X=9560000 $Y=3808000
X1923 24 1898 mux21_ni $T=9568000 1952000 0 0 $X=9568000 $Y=1952000
X1924 24 1899 mux21_ni $T=9584000 7520000 0 0 $X=9584000 $Y=7520000
X1925 24 1900 mux21_ni $T=9616000 9144000 0 0 $X=9616000 $Y=9144000
X1926 24 1901 mux21_ni $T=9624000 3576000 0 0 $X=9624000 $Y=3576000
X1927 24 1902 mux21_ni $T=9632000 1720000 0 0 $X=9632000 $Y=1720000
X1928 24 1903 mux21_ni $T=9656000 560000 0 0 $X=9656000 $Y=560000
X1929 24 1904 mux21_ni $T=9656000 3344000 0 0 $X=9656000 $Y=3344000
X1930 24 1905 mux21_ni $T=9664000 3112000 0 0 $X=9664000 $Y=3112000
X1931 24 1906 mux21_ni $T=9680000 10304000 0 0 $X=9680000 $Y=10304000
X1932 24 1907 mux21_ni $T=9696000 4736000 0 0 $X=9696000 $Y=4736000
X1933 24 1908 mux21_ni $T=9720000 10072000 0 0 $X=9720000 $Y=10072000
X1934 24 1909 mux21_ni $T=9728000 11232000 0 0 $X=9728000 $Y=11232000
X1935 24 1910 mux21_ni $T=9736000 7752000 0 0 $X=9736000 $Y=7752000
X1936 24 1911 mux21_ni $T=9784000 1488000 0 0 $X=9784000 $Y=1488000
X1937 24 1912 mux21_ni $T=9808000 96000 0 0 $X=9808000 $Y=96000
X1938 24 1913 mux21_ni $T=9808000 328000 0 0 $X=9808000 $Y=328000
X1939 24 1914 mux21_ni $T=9816000 2648000 0 0 $X=9816000 $Y=2648000
X1940 24 1915 mux21_ni $T=9816000 2880000 0 0 $X=9816000 $Y=2880000
X1941 24 1916 mux21_ni $T=9876000 7056000 1 180 $X=9816000 $Y=7056000
X1942 24 1917 mux21_ni $T=9824000 5896000 0 0 $X=9824000 $Y=5896000
X1943 24 1918 mux21_ni $T=9824000 6592000 0 0 $X=9824000 $Y=6592000
X1944 24 1919 mux21_ni $T=9824000 9840000 0 0 $X=9824000 $Y=9840000
X1945 24 1920 mux21_ni $T=9832000 8216000 0 0 $X=9832000 $Y=8216000
X1946 24 1921 mux21_ni $T=9840000 2416000 0 0 $X=9840000 $Y=2416000
X1947 24 1922 mux21_ni $T=9840000 10768000 0 0 $X=9840000 $Y=10768000
X1948 24 1923 mux21_ni $T=9908000 6128000 1 180 $X=9848000 $Y=6128000
X1949 24 1924 mux21_ni $T=9864000 3808000 0 0 $X=9864000 $Y=3808000
X1950 24 1925 mux21_ni $T=9864000 8680000 0 0 $X=9864000 $Y=8680000
X1951 24 1926 mux21_ni $T=9872000 1952000 0 0 $X=9872000 $Y=1952000
X1952 24 1927 mux21_ni $T=9872000 4272000 0 0 $X=9872000 $Y=4272000
X1953 24 1928 mux21_ni $T=9888000 6824000 0 0 $X=9888000 $Y=6824000
X1954 24 1929 mux21_ni $T=9888000 11928000 0 0 $X=9888000 $Y=11928000
X1955 24 1930 mux21_ni $T=9928000 3576000 0 0 $X=9928000 $Y=3576000
X1956 24 1931 mux21_ni $T=9988000 11000000 1 180 $X=9928000 $Y=11000000
X1957 24 1932 mux21_ni $T=9936000 3344000 0 0 $X=9936000 $Y=3344000
X1958 24 1933 mux21_ni $T=9936000 7056000 0 0 $X=9936000 $Y=7056000
X1959 24 1934 mux21_ni $T=9944000 6128000 0 0 $X=9944000 $Y=6128000
X1960 24 1935 mux21_ni $T=9952000 4504000 0 0 $X=9952000 $Y=4504000
X1961 24 1936 mux21_ni $T=9952000 11464000 0 0 $X=9952000 $Y=11464000
X1962 24 1937 mux21_ni $T=9960000 12392000 0 0 $X=9960000 $Y=12392000
X1963 24 1938 mux21_ni $T=9976000 3112000 0 0 $X=9976000 $Y=3112000
X1964 24 1939 mux21_ni $T=10024000 10072000 0 0 $X=10024000 $Y=10072000
X1965 24 1940 mux21_ni $T=10040000 4968000 0 0 $X=10040000 $Y=4968000
X1966 24 1941 mux21_ni $T=10112000 96000 0 0 $X=10112000 $Y=96000
X1967 24 1942 mux21_ni $T=10112000 12160000 0 0 $X=10112000 $Y=12160000
X1968 24 1943 mux21_ni $T=10120000 2880000 0 0 $X=10120000 $Y=2880000
X1969 24 1944 mux21_ni $T=10120000 10304000 0 0 $X=10120000 $Y=10304000
X1970 24 1945 mux21_ni $T=10136000 7288000 0 0 $X=10136000 $Y=7288000
X1971 24 1946 mux21_ni $T=10136000 7520000 0 0 $X=10136000 $Y=7520000
X1972 24 1947 mux21_ni $T=10144000 8680000 0 0 $X=10144000 $Y=8680000
X1973 24 1948 mux21_ni $T=10152000 9376000 0 0 $X=10152000 $Y=9376000
X1974 24 1949 mux21_ni $T=10228000 5432000 1 180 $X=10168000 $Y=5432000
X1975 24 1950 mux21_ni $T=10168000 6360000 0 0 $X=10168000 $Y=6360000
X1976 24 1951 mux21_ni $T=10168000 8912000 0 0 $X=10168000 $Y=8912000
X1977 24 1952 mux21_ni $T=10184000 2416000 0 0 $X=10184000 $Y=2416000
X1978 24 1953 mux21_ni $T=10248000 6128000 0 0 $X=10248000 $Y=6128000
X1979 24 1954 mux21_ni $T=10324000 7752000 1 180 $X=10264000 $Y=7752000
X1980 24 1955 mux21_ni $T=10332000 5664000 1 180 $X=10272000 $Y=5664000
X1981 24 1956 mux21_ni $T=10356000 11000000 1 180 $X=10296000 $Y=11000000
X1982 24 1957 mux21_ni $T=10380000 8216000 1 180 $X=10320000 $Y=8216000
X1983 24 1958 mux21_ni $T=10328000 7752000 0 0 $X=10328000 $Y=7752000
X1984 24 1959 mux21_ni $T=10388000 10072000 1 180 $X=10328000 $Y=10072000
X1985 24 1960 mux21_ni $T=10412000 13320000 1 180 $X=10352000 $Y=13320000
X1986 24 1961 mux21_ni $T=10360000 5896000 0 0 $X=10360000 $Y=5896000
X1987 24 1962 mux21_ni $T=10360000 8448000 0 0 $X=10360000 $Y=8448000
X1988 24 1963 mux21_ni $T=10360000 10536000 0 0 $X=10360000 $Y=10536000
X1989 24 1964 mux21_ni $T=10360000 11928000 0 0 $X=10360000 $Y=11928000
X1990 24 1965 mux21_ni $T=10384000 8216000 0 0 $X=10384000 $Y=8216000
X1991 24 1966 mux21_ni $T=10384000 9608000 0 0 $X=10384000 $Y=9608000
X1992 24 1967 mux21_ni $T=10400000 560000 0 0 $X=10400000 $Y=560000
X1993 24 1968 mux21_ni $T=10400000 12160000 0 0 $X=10400000 $Y=12160000
X1994 24 1969 mux21_ni $T=10416000 4504000 0 0 $X=10416000 $Y=4504000
X1995 24 1970 mux21_ni $T=10416000 13320000 0 0 $X=10416000 $Y=13320000
X1996 24 1971 mux21_ni $T=10424000 5896000 0 0 $X=10424000 $Y=5896000
X1997 24 1972 mux21_ni $T=10424000 9840000 0 0 $X=10424000 $Y=9840000
X1998 24 1973 mux21_ni $T=10484000 11464000 1 180 $X=10424000 $Y=11464000
X1999 24 1974 mux21_ni $T=10432000 12392000 0 0 $X=10432000 $Y=12392000
X2000 24 1975 mux21_ni $T=10440000 96000 0 0 $X=10440000 $Y=96000
X2001 24 1976 mux21_ni $T=10440000 6824000 0 0 $X=10440000 $Y=6824000
X2002 24 1977 mux21_ni $T=10448000 10768000 0 0 $X=10448000 $Y=10768000
X2003 24 1978 mux21_ni $T=10516000 3344000 1 180 $X=10456000 $Y=3344000
X2004 24 1979 mux21_ni $T=10456000 5200000 0 0 $X=10456000 $Y=5200000
X2005 24 1980 mux21_ni $T=10472000 8680000 0 0 $X=10472000 $Y=8680000
X2006 24 1981 mux21_ni $T=10540000 1720000 1 180 $X=10480000 $Y=1720000
X2007 24 1982 mux21_ni $T=10488000 2880000 0 0 $X=10488000 $Y=2880000
X2008 24 1983 mux21_ni $T=10488000 11000000 0 0 $X=10488000 $Y=11000000
X2009 24 1984 mux21_ni $T=10488000 12856000 0 0 $X=10488000 $Y=12856000
X2010 24 1985 mux21_ni $T=10496000 10072000 0 0 $X=10496000 $Y=10072000
X2011 24 1986 mux21_ni $T=10512000 5432000 0 0 $X=10512000 $Y=5432000
X2012 24 1987 mux21_ni $T=10520000 560000 0 0 $X=10520000 $Y=560000
X2013 24 1988 mux21_ni $T=10520000 2184000 0 0 $X=10520000 $Y=2184000
X2014 24 1989 mux21_ni $T=10536000 12624000 0 0 $X=10536000 $Y=12624000
X2015 24 1990 mux21_ni $T=10628000 792000 1 180 $X=10568000 $Y=792000
X2016 24 1991 mux21_ni $T=10628000 7984000 1 180 $X=10568000 $Y=7984000
X2017 24 1992 mux21_ni $T=10576000 3344000 0 0 $X=10576000 $Y=3344000
X2018 24 1993 mux21_ni $T=10584000 96000 0 0 $X=10584000 $Y=96000
X2019 24 1994 mux21_ni $T=10584000 560000 0 0 $X=10584000 $Y=560000
X2020 24 1995 mux21_ni $T=10584000 1024000 0 0 $X=10584000 $Y=1024000
X2021 24 1996 mux21_ni $T=10592000 4968000 0 0 $X=10592000 $Y=4968000
X2022 24 1997 mux21_ni $T=10632000 7520000 0 0 $X=10632000 $Y=7520000
X2023 24 1998 mux21_ni $T=10640000 3576000 0 0 $X=10640000 $Y=3576000
X2024 24 1999 mux21_ni $T=10648000 96000 0 0 $X=10648000 $Y=96000
X2025 24 2000 mux21_ni $T=10648000 4272000 0 0 $X=10648000 $Y=4272000
X2026 24 2001 mux21_ni $T=10680000 4040000 0 0 $X=10680000 $Y=4040000
X2027 24 2002 mux21_ni $T=10680000 6592000 0 0 $X=10680000 $Y=6592000
X2028 24 2003 mux21_ni $T=10688000 7288000 0 0 $X=10688000 $Y=7288000
X2029 24 2004 mux21_ni $T=10712000 6360000 0 0 $X=10712000 $Y=6360000
X2030 24 2005 mux21_ni $T=10744000 4040000 0 0 $X=10744000 $Y=4040000
X2031 24 2006 mux21_ni $T=10744000 4736000 0 0 $X=10744000 $Y=4736000
X2032 24 2007 mux21_ni $T=10804000 8216000 1 180 $X=10744000 $Y=8216000
X2033 24 2008 mux21_ni $T=10760000 3576000 0 0 $X=10760000 $Y=3576000
X2034 24 2009 mux21_ni $T=10768000 9840000 0 0 $X=10768000 $Y=9840000
X2035 24 2010 mux21_ni $T=10768000 11232000 0 0 $X=10768000 $Y=11232000
X2036 24 2011 mux21_ni $T=10784000 10536000 0 0 $X=10784000 $Y=10536000
X2037 24 2012 mux21_ni $T=10792000 96000 0 0 $X=10792000 $Y=96000
X2038 24 2013 mux21_ni $T=10792000 9608000 0 0 $X=10792000 $Y=9608000
X2039 24 2014 mux21_ni $T=10816000 5432000 0 0 $X=10816000 $Y=5432000
X2040 24 2015 mux21_ni $T=10832000 3112000 0 0 $X=10832000 $Y=3112000
X2041 24 2016 mux21_ni $T=10892000 13320000 1 180 $X=10832000 $Y=13320000
X2042 24 2017 mux21_ni $T=10848000 7056000 0 0 $X=10848000 $Y=7056000
X2043 24 2018 mux21_ni $T=10848000 7984000 0 0 $X=10848000 $Y=7984000
X2044 24 2019 mux21_ni $T=10916000 96000 1 180 $X=10856000 $Y=96000
X2045 24 2020 mux21_ni $T=10856000 10304000 0 0 $X=10856000 $Y=10304000
X2046 24 2021 mux21_ni $T=10856000 10768000 0 0 $X=10856000 $Y=10768000
X2047 24 2022 mux21_ni $T=10864000 7752000 0 0 $X=10864000 $Y=7752000
X2048 24 2023 mux21_ni $T=10924000 11696000 1 180 $X=10864000 $Y=11696000
X2049 24 2024 mux21_ni $T=10872000 5200000 0 0 $X=10872000 $Y=5200000
X2050 24 2025 mux21_ni $T=10880000 10072000 0 0 $X=10880000 $Y=10072000
X2051 24 2026 mux21_ni $T=10888000 4504000 0 0 $X=10888000 $Y=4504000
X2052 24 2027 mux21_ni $T=10912000 6128000 0 0 $X=10912000 $Y=6128000
X2053 24 2028 mux21_ni $T=10912000 7056000 0 0 $X=10912000 $Y=7056000
X2054 24 2029 mux21_ni $T=10928000 9144000 0 0 $X=10928000 $Y=9144000
X2055 24 2030 mux21_ni $T=10928000 13320000 0 0 $X=10928000 $Y=13320000
X2056 24 2031 mux21_ni $T=10936000 5664000 0 0 $X=10936000 $Y=5664000
X2057 24 2032 mux21_ni $T=10944000 8912000 0 0 $X=10944000 $Y=8912000
X2058 24 2033 mux21_ni $T=10944000 11000000 0 0 $X=10944000 $Y=11000000
X2059 24 2034 mux21_ni $T=11020000 96000 1 180 $X=10960000 $Y=96000
X2060 24 2035 mux21_ni $T=10976000 2648000 0 0 $X=10976000 $Y=2648000
X2061 24 2036 mux21_ni $T=10984000 6592000 0 0 $X=10984000 $Y=6592000
X2062 24 2037 mux21_ni $T=10992000 7288000 0 0 $X=10992000 $Y=7288000
X2063 24 2038 mux21_ni $T=10992000 7520000 0 0 $X=10992000 $Y=7520000
X2064 24 2039 mux21_ni $T=11000000 5664000 0 0 $X=11000000 $Y=5664000
X2065 24 2040 mux21_ni $T=11016000 12856000 0 0 $X=11016000 $Y=12856000
X2066 24 2041 mux21_ni $T=11024000 8680000 0 0 $X=11024000 $Y=8680000
X2067 24 2042 mux21_ni $T=11100000 1720000 1 180 $X=11040000 $Y=1720000
X2068 24 2043 mux21_ni $T=11048000 2880000 0 0 $X=11048000 $Y=2880000
X2069 24 2044 mux21_ni $T=11048000 4040000 0 0 $X=11048000 $Y=4040000
X2070 24 2045 mux21_ni $T=11056000 328000 0 0 $X=11056000 $Y=328000
X2071 24 2046 mux21_ni $T=11124000 96000 1 180 $X=11064000 $Y=96000
X2072 24 2047 mux21_ni $T=11072000 1024000 0 0 $X=11072000 $Y=1024000
X2073 24 2048 mux21_ni $T=11148000 8216000 1 180 $X=11088000 $Y=8216000
X2074 24 2049 mux21_ni $T=11088000 12160000 0 0 $X=11088000 $Y=12160000
X2075 24 2050 mux21_ni $T=11096000 1256000 0 0 $X=11096000 $Y=1256000
X2076 24 2051 mux21_ni $T=11104000 11232000 0 0 $X=11104000 $Y=11232000
X2077 24 2052 mux21_ni $T=11188000 96000 1 180 $X=11128000 $Y=96000
X2078 24 2053 mux21_ni $T=11136000 1720000 0 0 $X=11136000 $Y=1720000
X2079 24 2054 mux21_ni $T=11152000 8216000 0 0 $X=11152000 $Y=8216000
X2080 24 2055 mux21_ni $T=11152000 12392000 0 0 $X=11152000 $Y=12392000
X2081 24 2056 mux21_ni $T=11220000 11696000 1 180 $X=11160000 $Y=11696000
X2082 24 2057 mux21_ni $T=11236000 2416000 1 180 $X=11176000 $Y=2416000
X2083 24 2058 mux21_ni $T=11176000 3112000 0 0 $X=11176000 $Y=3112000
X2084 24 2059 mux21_ni $T=11176000 5432000 0 0 $X=11176000 $Y=5432000
X2085 24 2060 mux21_ni $T=11200000 1256000 0 0 $X=11200000 $Y=1256000
X2086 24 2061 mux21_ni $T=11216000 7056000 0 0 $X=11216000 $Y=7056000
X2087 24 2062 mux21_ni $T=11224000 8448000 0 0 $X=11224000 $Y=8448000
X2088 24 2063 mux21_ni $T=11224000 11696000 0 0 $X=11224000 $Y=11696000
X2089 24 2064 mux21_ni $T=11240000 3112000 0 0 $X=11240000 $Y=3112000
X2090 24 2065 mux21_ni $T=11240000 4272000 0 0 $X=11240000 $Y=4272000
X2091 24 2066 mux21_ni $T=11248000 8912000 0 0 $X=11248000 $Y=8912000
X2092 24 2067 mux21_ni $T=11256000 6128000 0 0 $X=11256000 $Y=6128000
X2093 24 2068 mux21_ni $T=11304000 328000 0 0 $X=11304000 $Y=328000
X2094 24 2069 mux21_ni $T=11304000 1256000 0 0 $X=11304000 $Y=1256000
X2095 24 2070 mux21_ni $T=11304000 6360000 0 0 $X=11304000 $Y=6360000
X2096 24 2071 mux21_ni $T=11336000 4968000 0 0 $X=11336000 $Y=4968000
X2097 24 2072 mux21_ni $T=11344000 1024000 0 0 $X=11344000 $Y=1024000
X2098 24 2073 mux21_ni $T=11352000 96000 0 0 $X=11352000 $Y=96000
X2099 24 2074 mux21_ni $T=11420000 4040000 1 180 $X=11360000 $Y=4040000
X2100 24 2075 mux21_ni $T=11428000 13320000 1 180 $X=11368000 $Y=13320000
X2101 24 2076 mux21_ni $T=11384000 560000 0 0 $X=11384000 $Y=560000
X2102 24 2077 mux21_ni $T=11384000 4504000 0 0 $X=11384000 $Y=4504000
X2103 24 2078 mux21_ni $T=11408000 328000 0 0 $X=11408000 $Y=328000
X2104 24 2079 mux21_ni $T=11408000 1024000 0 0 $X=11408000 $Y=1024000
X2105 24 2080 mux21_ni $T=11408000 10304000 0 0 $X=11408000 $Y=10304000
X2106 24 2081 mux21_ni $T=11416000 792000 0 0 $X=11416000 $Y=792000
X2107 24 2082 mux21_ni $T=11424000 2184000 0 0 $X=11424000 $Y=2184000
X2108 24 2083 mux21_ni $T=11424000 4040000 0 0 $X=11424000 $Y=4040000
X2109 24 2084 mux21_ni $T=11484000 6592000 1 180 $X=11424000 $Y=6592000
X2110 24 2085 mux21_ni $T=11492000 1256000 1 180 $X=11432000 $Y=1256000
X2111 24 2086 mux21_ni $T=11492000 3576000 1 180 $X=11432000 $Y=3576000
X2112 24 2087 mux21_ni $T=11492000 7984000 1 180 $X=11432000 $Y=7984000
X2113 24 2088 mux21_ni $T=11448000 560000 0 0 $X=11448000 $Y=560000
X2114 24 2089 mux21_ni $T=11516000 12392000 1 180 $X=11456000 $Y=12392000
X2115 24 2090 mux21_ni $T=11472000 328000 0 0 $X=11472000 $Y=328000
X2116 24 2091 mux21_ni $T=11472000 1024000 0 0 $X=11472000 $Y=1024000
X2117 24 2092 mux21_ni $T=11488000 11464000 0 0 $X=11488000 $Y=11464000
X2118 24 2093 mux21_ni $T=11496000 96000 0 0 $X=11496000 $Y=96000
X2119 24 2094 mux21_ni $T=11556000 1256000 1 180 $X=11496000 $Y=1256000
X2120 24 2095 mux21_ni $T=11496000 9840000 0 0 $X=11496000 $Y=9840000
X2121 24 2096 mux21_ni $T=11588000 7056000 1 180 $X=11528000 $Y=7056000
X2122 24 2097 mux21_ni $T=11528000 9608000 0 0 $X=11528000 $Y=9608000
X2123 24 2098 mux21_ni $T=11536000 328000 0 0 $X=11536000 $Y=328000
X2124 24 2099 mux21_ni $T=11536000 5200000 0 0 $X=11536000 $Y=5200000
X2125 24 2100 mux21_ni $T=11604000 792000 1 180 $X=11544000 $Y=792000
X2126 24 2101 mux21_ni $T=11544000 7288000 0 0 $X=11544000 $Y=7288000
X2127 24 2102 mux21_ni $T=11612000 560000 1 180 $X=11552000 $Y=560000
X2128 24 2103 mux21_ni $T=11552000 4272000 0 0 $X=11552000 $Y=4272000
X2129 24 2104 mux21_ni $T=11552000 8912000 0 0 $X=11552000 $Y=8912000
X2130 24 2105 mux21_ni $T=11620000 2648000 1 180 $X=11560000 $Y=2648000
X2131 24 2106 mux21_ni $T=11600000 328000 0 0 $X=11600000 $Y=328000
X2132 24 2107 mux21_ni $T=11660000 1256000 1 180 $X=11600000 $Y=1256000
X2133 24 2108 mux21_ni $T=11600000 11232000 0 0 $X=11600000 $Y=11232000
X2134 24 2109 mux21_ni $T=11616000 8912000 0 0 $X=11616000 $Y=8912000
X2135 24 2110 mux21_ni $T=11640000 13088000 0 0 $X=11640000 $Y=13088000
X2136 24 2111 mux21_ni $T=11708000 792000 1 180 $X=11648000 $Y=792000
X2137 24 2112 mux21_ni $T=11664000 4968000 0 0 $X=11664000 $Y=4968000
X2138 24 2113 mux21_ni $T=11664000 6360000 0 0 $X=11664000 $Y=6360000
X2139 24 2114 mux21_ni $T=11664000 11000000 0 0 $X=11664000 $Y=11000000
X2140 24 2115 mux21_ni $T=11680000 96000 0 0 $X=11680000 $Y=96000
X2141 24 2116 mux21_ni $T=11680000 3808000 0 0 $X=11680000 $Y=3808000
X2142 24 2117 mux21_ni $T=11680000 8912000 0 0 $X=11680000 $Y=8912000
X2143 24 2118 mux21_ni $T=11756000 7752000 1 180 $X=11696000 $Y=7752000
X2144 24 2119 mux21_ni $T=11696000 11696000 0 0 $X=11696000 $Y=11696000
X2145 24 2120 mux21_ni $T=11704000 13320000 0 0 $X=11704000 $Y=13320000
X2146 24 2121 mux21_ni $T=11712000 2648000 0 0 $X=11712000 $Y=2648000
X2147 24 2122 mux21_ni $T=11720000 8448000 0 0 $X=11720000 $Y=8448000
X2148 24 2123 mux21_ni $T=11780000 10304000 1 180 $X=11720000 $Y=10304000
X2149 24 2124 mux21_ni $T=11720000 10768000 0 0 $X=11720000 $Y=10768000
X2150 24 2125 mux21_ni $T=11728000 1952000 0 0 $X=11728000 $Y=1952000
X2151 24 2126 mux21_ni $T=11728000 2416000 0 0 $X=11728000 $Y=2416000
X2152 24 2127 mux21_ni $T=11728000 4968000 0 0 $X=11728000 $Y=4968000
X2153 24 2128 mux21_ni $T=11728000 12392000 0 0 $X=11728000 $Y=12392000
X2154 24 2129 mux21_ni $T=11804000 96000 1 180 $X=11744000 $Y=96000
X2155 24 2130 mux21_ni $T=11744000 5896000 0 0 $X=11744000 $Y=5896000
X2156 24 2131 mux21_ni $T=11760000 2880000 0 0 $X=11760000 $Y=2880000
X2157 24 2132 mux21_ni $T=11768000 12624000 0 0 $X=11768000 $Y=12624000
X2158 24 2133 mux21_ni $T=11768000 13552000 0 0 $X=11768000 $Y=13552000
X2159 24 2134 mux21_ni $T=11784000 4040000 0 0 $X=11784000 $Y=4040000
X2160 24 2135 mux21_ni $T=11792000 7520000 0 0 $X=11792000 $Y=7520000
X2161 24 2136 mux21_ni $T=11800000 3344000 0 0 $X=11800000 $Y=3344000
X2162 24 2137 mux21_ni $T=11800000 3576000 0 0 $X=11800000 $Y=3576000
X2163 24 2138 mux21_ni $T=11808000 1720000 0 0 $X=11808000 $Y=1720000
X2164 24 2139 mux21_ni $T=11832000 792000 0 0 $X=11832000 $Y=792000
X2165 24 2140 mux21_ni $T=11832000 6824000 0 0 $X=11832000 $Y=6824000
X2166 24 2141 mux21_ni $T=11908000 96000 1 180 $X=11848000 $Y=96000
X2167 24 2142 mux21_ni $T=11856000 4272000 0 0 $X=11856000 $Y=4272000
X2168 24 2143 mux21_ni $T=11856000 7520000 0 0 $X=11856000 $Y=7520000
X2169 24 2144 mux21_ni $T=11864000 3344000 0 0 $X=11864000 $Y=3344000
X2170 24 2145 mux21_ni $T=11948000 1024000 1 180 $X=11888000 $Y=1024000
X2171 24 2146 mux21_ni $T=11896000 792000 0 0 $X=11896000 $Y=792000
X2172 24 2147 mux21_ni $T=11928000 13088000 0 0 $X=11928000 $Y=13088000
X2173 24 2148 mux21_ni $T=11944000 328000 0 0 $X=11944000 $Y=328000
X2174 24 2149 mux21_ni $T=11944000 8680000 0 0 $X=11944000 $Y=8680000
X2175 24 2150 mux21_ni $T=11968000 6592000 0 0 $X=11968000 $Y=6592000
X2176 24 2151 mux21_ni $T=12036000 560000 1 180 $X=11976000 $Y=560000
X2177 24 2152 mux21_ni $T=11984000 1256000 0 0 $X=11984000 $Y=1256000
X2178 24 2153 mux21_ni $T=11984000 12160000 0 0 $X=11984000 $Y=12160000
X2179 24 2154 mux21_ni $T=11992000 96000 0 0 $X=11992000 $Y=96000
X2180 24 2155 mux21_ni $T=12000000 792000 0 0 $X=12000000 $Y=792000
X2181 24 2156 mux21_ni $T=12008000 328000 0 0 $X=12008000 $Y=328000
X2182 24 2157 mux21_ni $T=12068000 8680000 1 180 $X=12008000 $Y=8680000
X2183 24 2158 mux21_ni $T=12032000 2184000 0 0 $X=12032000 $Y=2184000
X2184 24 2159 mux21_ni $T=12032000 2416000 0 0 $X=12032000 $Y=2416000
X2185 24 2160 mux21_ni $T=12032000 7056000 0 0 $X=12032000 $Y=7056000
X2186 24 2161 mux21_ni $T=12032000 11696000 0 0 $X=12032000 $Y=11696000
X2187 24 2162 mux21_ni $T=12032000 12856000 0 0 $X=12032000 $Y=12856000
X2188 24 2163 mux21_ni $T=12040000 3808000 0 0 $X=12040000 $Y=3808000
X2189 24 2164 mux21_ni $T=12048000 7288000 0 0 $X=12048000 $Y=7288000
X2190 24 2165 mux21_ni $T=12156000 2880000 1 180 $X=12096000 $Y=2880000
X2191 24 2166 mux21_ni $T=12096000 6824000 0 0 $X=12096000 $Y=6824000
X2192 24 2167 mux21_ni $T=12096000 13552000 0 0 $X=12096000 $Y=13552000
X2193 24 2168 mux21_ni $T=12104000 3808000 0 0 $X=12104000 $Y=3808000
X2194 24 2169 mux21_ni $T=12104000 13088000 0 0 $X=12104000 $Y=13088000
X2195 24 2170 mux21_ni $T=12172000 1256000 1 180 $X=12112000 $Y=1256000
X2196 24 2171 mux21_ni $T=12172000 8680000 1 180 $X=12112000 $Y=8680000
X2197 24 2172 mux21_ni $T=12128000 1720000 0 0 $X=12128000 $Y=1720000
X2198 24 2173 mux21_ni $T=12136000 7056000 0 0 $X=12136000 $Y=7056000
X2199 24 2174 mux21_ni $T=12136000 12624000 0 0 $X=12136000 $Y=12624000
X2200 24 2175 mux21_ni $T=12168000 3344000 0 0 $X=12168000 $Y=3344000
X2201 24 2176 mux21_ni $T=12176000 328000 0 0 $X=12176000 $Y=328000
X2202 24 2177 mux21_ni $T=12236000 7288000 1 180 $X=12176000 $Y=7288000
X2203 24 2178 mux21_ni $T=12200000 12624000 0 0 $X=12200000 $Y=12624000
X2204 24 2179 mux21_ni $T=12208000 13088000 0 0 $X=12208000 $Y=13088000
X2205 24 2180 mux21_ni $T=12216000 96000 0 0 $X=12216000 $Y=96000
X2206 24 2181 mux21_ni $T=12276000 1256000 1 180 $X=12216000 $Y=1256000
X2207 24 2182 mux21_ni $T=12216000 4272000 0 0 $X=12216000 $Y=4272000
X2208 24 2183 mux21_ni $T=12276000 7520000 1 180 $X=12216000 $Y=7520000
X2209 24 2184 mux21_ni $T=12216000 8448000 0 0 $X=12216000 $Y=8448000
X2210 24 2185 mux21_ni $T=12216000 8912000 0 0 $X=12216000 $Y=8912000
X2211 24 2186 mux21_ni $T=12216000 10768000 0 0 $X=12216000 $Y=10768000
X2212 24 2187 mux21_ni $T=12216000 11928000 0 0 $X=12216000 $Y=11928000
X2213 24 2188 mux21_ni $T=12224000 1952000 0 0 $X=12224000 $Y=1952000
X2214 24 2189 mux21_ni $T=12224000 11000000 0 0 $X=12224000 $Y=11000000
X2215 24 2190 mux21_ni $T=12232000 3344000 0 0 $X=12232000 $Y=3344000
X2216 24 2191 mux21_ni $T=12240000 328000 0 0 $X=12240000 $Y=328000
X2217 24 2192 mux21_ni $T=12300000 560000 1 180 $X=12240000 $Y=560000
X2218 24 2193 mux21_ni $T=12240000 792000 0 0 $X=12240000 $Y=792000
X2219 24 2194 mux21_ni $T=12324000 7056000 1 180 $X=12264000 $Y=7056000
X2220 24 2195 mux21_ni $T=12264000 10072000 0 0 $X=12264000 $Y=10072000
X2221 24 2196 mux21_ni $T=12264000 11232000 0 0 $X=12264000 $Y=11232000
X2222 24 2197 mux21_ni $T=12264000 12392000 0 0 $X=12264000 $Y=12392000
X2223 24 2198 mux21_ni $T=12332000 5664000 1 180 $X=12272000 $Y=5664000
X2224 24 2199 mux21_ni $T=12272000 5896000 0 0 $X=12272000 $Y=5896000
X2225 24 2200 mux21_ni $T=12272000 13088000 0 0 $X=12272000 $Y=13088000
X2226 24 2201 mux21_ni $T=12340000 96000 1 180 $X=12280000 $Y=96000
X2227 24 2202 mux21_ni $T=12280000 2648000 0 0 $X=12280000 $Y=2648000
X2228 24 2203 mux21_ni $T=12280000 3808000 0 0 $X=12280000 $Y=3808000
X2229 24 2204 mux21_ni $T=12280000 4272000 0 0 $X=12280000 $Y=4272000
X2230 24 2205 mux21_ni $T=12280000 4736000 0 0 $X=12280000 $Y=4736000
X2231 24 2206 mux21_ni $T=12280000 4968000 0 0 $X=12280000 $Y=4968000
X2232 24 2207 mux21_ni $T=12280000 5200000 0 0 $X=12280000 $Y=5200000
X2233 24 2208 mux21_ni $T=12280000 6128000 0 0 $X=12280000 $Y=6128000
X2234 24 2209 mux21_ni $T=12280000 6592000 0 0 $X=12280000 $Y=6592000
X2235 24 2210 mux21_ni $T=12340000 7288000 1 180 $X=12280000 $Y=7288000
X2236 24 2211 mux21_ni $T=12280000 7752000 0 0 $X=12280000 $Y=7752000
X2237 24 2212 mux21_ni $T=12280000 7984000 0 0 $X=12280000 $Y=7984000
X2238 24 2213 mux21_ni $T=12280000 8448000 0 0 $X=12280000 $Y=8448000
X2239 24 2214 mux21_ni $T=12280000 8912000 0 0 $X=12280000 $Y=8912000
X2240 24 2215 mux21_ni $T=12280000 9376000 0 0 $X=12280000 $Y=9376000
X2241 24 2216 mux21_ni $T=12280000 9608000 0 0 $X=12280000 $Y=9608000
X2242 24 2217 mux21_ni $T=12280000 9840000 0 0 $X=12280000 $Y=9840000
X2243 24 2218 mux21_ni $T=12280000 10304000 0 0 $X=12280000 $Y=10304000
X2244 24 2219 mux21_ni $T=12280000 10768000 0 0 $X=12280000 $Y=10768000
X2245 24 2220 mux21_ni $T=12280000 11928000 0 0 $X=12280000 $Y=11928000
X2246 24 2221 mux21_ni $T=12280000 12160000 0 0 $X=12280000 $Y=12160000
X2247 24 2222 mux21_ni $T=12348000 1024000 1 180 $X=12288000 $Y=1024000
X2248 24 2223 mux21_ni $T=12380000 1256000 1 180 $X=12320000 $Y=1256000
X2249 24 2224 mux21_ni $T=12380000 7520000 1 180 $X=12320000 $Y=7520000
X2250 24 2225 mux21_ni $T=12388000 7056000 1 180 $X=12328000 $Y=7056000
X2251 24 2226 mux21_ni $T=12336000 5896000 0 0 $X=12336000 $Y=5896000
X2252 24 2227 mux21_ni $T=12412000 1024000 1 180 $X=12352000 $Y=1024000
X2253 24 2228 mux21_ni $T=12420000 1488000 1 180 $X=12360000 $Y=1488000
X2254 24 2229 mux21_ni $T=12444000 96000 1 180 $X=12384000 $Y=96000
X2255 24 2230 mux21_ni $T=12444000 328000 1 180 $X=12384000 $Y=328000
X2256 24 2231 mux21_ni $T=12444000 1256000 1 180 $X=12384000 $Y=1256000
X2257 24 2232 mux21_ni $T=12444000 6824000 1 180 $X=12384000 $Y=6824000
X2258 24 2233 mux21_ni $T=12444000 7520000 1 180 $X=12384000 $Y=7520000
X2259 24 2234 mux21_ni $T=12444000 8912000 1 180 $X=12384000 $Y=8912000
X2260 24 2235 mux21_ni $T=12484000 7056000 1 180 $X=12424000 $Y=7056000
X2261 24 2236 mux21_ni $T=12484000 7288000 1 180 $X=12424000 $Y=7288000
X2262 24 2237 mux21_ni $T=12484000 8680000 1 180 $X=12424000 $Y=8680000
X2263 24 2238 mux21 $T=152000 2648000 0 0 $X=152000 $Y=2648000
X2264 24 2239 mux21 $T=216000 2648000 0 0 $X=216000 $Y=2648000
X2265 24 2240 mux21 $T=500500 2880000 1 180 $X=440000 $Y=2880000
X2266 24 2241 mux21 $T=568000 1024000 0 0 $X=568000 $Y=1024000
X2267 24 2242 mux21 $T=740500 2184000 1 180 $X=680000 $Y=2184000
X2268 24 2243 mux21 $T=912000 792000 0 0 $X=912000 $Y=792000
X2269 24 2244 mux21 $T=1144000 328000 0 0 $X=1144000 $Y=328000
X2270 24 2245 mux21 $T=1340500 3344000 1 180 $X=1280000 $Y=3344000
X2271 24 2246 mux21 $T=1432000 2184000 0 0 $X=1432000 $Y=2184000
X2272 24 2247 mux21 $T=1488000 2416000 0 0 $X=1488000 $Y=2416000
X2273 24 2248 mux21 $T=1568000 1952000 0 0 $X=1568000 $Y=1952000
X2274 24 2249 mux21 $T=1608000 1256000 0 0 $X=1608000 $Y=1256000
X2275 24 2250 mux21 $T=1880000 1488000 0 0 $X=1880000 $Y=1488000
X2276 24 2251 mux21 $T=1968000 1024000 0 0 $X=1968000 $Y=1024000
X2277 24 2252 mux21 $T=2440000 1488000 0 0 $X=2440000 $Y=1488000
X2278 24 2253 mux21 $T=2548500 1952000 1 180 $X=2488000 $Y=1952000
X2279 24 2254 mux21 $T=2564500 1488000 1 180 $X=2504000 $Y=1488000
X2280 24 2255 mux21 $T=2652500 3112000 1 180 $X=2592000 $Y=3112000
X2281 24 2256 mux21 $T=2720000 1256000 0 0 $X=2720000 $Y=1256000
X2282 24 2257 mux21 $T=2860500 1024000 1 180 $X=2800000 $Y=1024000
X2283 24 2258 mux21 $T=2916500 328000 1 180 $X=2856000 $Y=328000
X2284 24 2259 mux21 $T=2972500 2184000 1 180 $X=2912000 $Y=2184000
X2285 24 2260 mux21 $T=2980500 328000 1 180 $X=2920000 $Y=328000
X2286 24 2261 mux21 $T=3100500 1952000 1 180 $X=3040000 $Y=1952000
X2287 24 2262 mux21 $T=3200000 328000 0 0 $X=3200000 $Y=328000
X2288 24 2263 mux21 $T=3488000 328000 0 0 $X=3488000 $Y=328000
X2289 24 2264 mux21 $T=3828500 328000 1 180 $X=3768000 $Y=328000
X2290 24 2265 mux21 $T=4164500 560000 1 180 $X=4104000 $Y=560000
X2291 24 2266 mux21 $T=4268500 328000 1 180 $X=4208000 $Y=328000
X2292 24 2267 mux21 $T=10528000 328000 0 0 $X=10528000 $Y=328000
X2293 24 2268 mux21 $T=10816000 328000 0 0 $X=10816000 $Y=328000
X2294 24 2269 mux21 $T=10840000 792000 0 0 $X=10840000 $Y=792000
X2295 24 2270 mux21 $T=10960000 792000 0 0 $X=10960000 $Y=792000
X2296 24 2271 mux21 $T=11192000 792000 0 0 $X=11192000 $Y=792000
X2297 24 2272 mux21 $T=11200000 328000 0 0 $X=11200000 $Y=328000
X2298 24 2273 mux21 $T=11360000 1720000 0 0 $X=11360000 $Y=1720000
X2299 24 2274 mux21 $T=11428500 1256000 1 180 $X=11368000 $Y=1256000
X2300 24 2275 mux21 $T=11540500 792000 1 180 $X=11480000 $Y=792000
X2301 24 2276 mux21 $T=11664000 328000 0 0 $X=11664000 $Y=328000
X2302 24 2277 mux21 $T=11848000 1488000 0 0 $X=11848000 $Y=1488000
X2303 24 2278 mux21 $T=12108500 1256000 1 180 $X=12048000 $Y=1256000
X2304 24 2279 mux21 $T=12132500 328000 1 180 $X=12072000 $Y=328000
X2305 24 2280 mux21 $T=12172500 7288000 1 180 $X=12112000 $Y=7288000
X2306 24 2281 mux21 $T=12184000 1024000 0 0 $X=12184000 $Y=1024000
X2307 24 2282 mux21 $T=12200000 7056000 0 0 $X=12200000 $Y=7056000
X2308 24 2283 mux21 $T=12444500 792000 1 180 $X=12384000 $Y=792000
X2309 24 2284 mux21 $T=12484500 560000 1 180 $X=12424000 $Y=560000
X2310 24 2285 mux21 $T=12484500 1488000 1 180 $X=12424000 $Y=1488000
X2311 24 2286 dffr $T=152000 5664000 0 0 $X=152000 $Y=5664000
X2312 24 2287 dffr $T=152000 6360000 0 0 $X=152000 $Y=6360000
X2313 24 2288 dffr $T=152000 13552000 0 0 $X=152000 $Y=13552000
X2314 24 2289 dffr $T=584000 9144000 1 180 $X=400000 $Y=9144000
X2315 24 2290 dffr $T=584000 9376000 1 180 $X=400000 $Y=9376000
X2316 24 2291 dffr $T=528000 4504000 0 0 $X=528000 $Y=4504000
X2317 24 2292 dffr $T=528000 4736000 0 0 $X=528000 $Y=4736000
X2318 24 2293 dffr $T=784000 9608000 1 180 $X=600000 $Y=9608000
X2319 24 2294 dffr $T=832000 6592000 1 180 $X=648000 $Y=6592000
X2320 24 2295 dffr $T=944000 8216000 1 180 $X=760000 $Y=8216000
X2321 24 2296 dffr $T=840000 4272000 0 0 $X=840000 $Y=4272000
X2322 24 2297 dffr $T=976000 5432000 0 0 $X=976000 $Y=5432000
X2323 24 2298 dffr $T=992000 13552000 0 0 $X=992000 $Y=13552000
X2324 24 2299 dffr $T=1032000 10304000 0 0 $X=1032000 $Y=10304000
X2325 24 2300 dffr $T=1192000 12624000 0 0 $X=1192000 $Y=12624000
X2326 24 2301 dffr $T=1440000 11000000 0 0 $X=1440000 $Y=11000000
X2327 24 2302 dffr $T=1496000 7056000 0 0 $X=1496000 $Y=7056000
X2328 24 2303 dffr $T=1672000 7752000 0 0 $X=1672000 $Y=7752000
X2329 24 2304 dffr $T=2368000 3576000 1 180 $X=2184000 $Y=3576000
X2330 24 2305 dffr $T=2416000 4968000 0 0 $X=2416000 $Y=4968000
X2331 24 2306 dffr $T=2456000 6592000 0 0 $X=2456000 $Y=6592000
X2332 24 2307 dffr $T=2472000 6128000 0 0 $X=2472000 $Y=6128000
X2333 24 2308 dffr $T=2704000 5664000 1 180 $X=2520000 $Y=5664000
X2334 24 2309 dffr $T=2816000 4504000 1 180 $X=2632000 $Y=4504000
X2335 24 2310 dffr $T=2648000 5200000 0 0 $X=2648000 $Y=5200000
X2336 24 2311 dffr $T=3000000 5664000 1 180 $X=2816000 $Y=5664000
X2337 24 2312 dffr $T=2856000 3808000 0 0 $X=2856000 $Y=3808000
X2338 24 2313 dffr $T=3184000 2880000 0 0 $X=3184000 $Y=2880000
X2339 24 2314 dffr $T=3464000 2880000 0 0 $X=3464000 $Y=2880000
X2340 24 2315 dffr $T=3520000 7984000 0 0 $X=3520000 $Y=7984000
X2341 24 2316 dffr $T=3864000 13088000 0 0 $X=3864000 $Y=13088000
X2342 24 168 dffr $T=3896000 328000 0 0 $X=3896000 $Y=328000
X2343 24 2317 dffr $T=3904000 4968000 0 0 $X=3904000 $Y=4968000
X2344 24 2318 dffr $T=4008000 1024000 0 0 $X=4008000 $Y=1024000
X2345 24 2319 dffr $T=4512000 1720000 0 0 $X=4512000 $Y=1720000
X2346 24 2320 dffr $T=4576000 10768000 0 0 $X=4576000 $Y=10768000
X2347 24 2321 dffr $T=4768000 6592000 1 180 $X=4584000 $Y=6592000
X2348 24 2322 dffr $T=5400000 792000 1 180 $X=5216000 $Y=792000
X2349 24 2323 dffr $T=5448000 328000 1 180 $X=5264000 $Y=328000
X2350 24 2324 dffr $T=5576000 11928000 1 180 $X=5392000 $Y=11928000
X2351 24 2325 dffr $T=5512000 96000 0 0 $X=5512000 $Y=96000
X2352 24 2326 dffr $T=6208000 96000 1 180 $X=6024000 $Y=96000
X2353 24 2327 dffr $T=6104000 11464000 0 0 $X=6104000 $Y=11464000
X2354 24 2328 dffr $T=6296000 10072000 1 180 $X=6112000 $Y=10072000
X2355 24 2329 dffr $T=6144000 792000 0 0 $X=6144000 $Y=792000
X2356 24 2330 dffr $T=6144000 11232000 0 0 $X=6144000 $Y=11232000
X2357 24 2331 dffr $T=6144000 11696000 0 0 $X=6144000 $Y=11696000
X2358 24 2332 dffr $T=6376000 4504000 1 180 $X=6192000 $Y=4504000
X2359 24 2333 dffr $T=6400000 7056000 0 0 $X=6400000 $Y=7056000
X2360 24 2334 dffr $T=6400000 8448000 0 0 $X=6400000 $Y=8448000
X2361 24 2335 dffr $T=6480000 2416000 0 0 $X=6480000 $Y=2416000
X2362 24 2336 dffr $T=6592000 8448000 0 0 $X=6592000 $Y=8448000
X2363 24 2337 dffr $T=6640000 5664000 0 0 $X=6640000 $Y=5664000
X2364 24 2338 dffr $T=6656000 11232000 0 0 $X=6656000 $Y=11232000
X2365 24 2339 dffr $T=6840000 12392000 0 0 $X=6840000 $Y=12392000
X2366 24 2340 dffr $T=6960000 8216000 0 0 $X=6960000 $Y=8216000
X2367 24 2341 dffr $T=7368000 13552000 0 0 $X=7368000 $Y=13552000
X2368 24 2342 dffr $T=7488000 96000 0 0 $X=7488000 $Y=96000
X2369 24 2343 dffr $T=7728000 3344000 1 180 $X=7544000 $Y=3344000
X2370 24 2344 dffr $T=8736000 4736000 1 180 $X=8552000 $Y=4736000
X2371 24 2345 dffr $T=8872000 12160000 0 0 $X=8872000 $Y=12160000
X2372 24 2346 dffr $T=9152000 3808000 1 180 $X=8968000 $Y=3808000
X2373 24 2347 dffr $T=9272000 4968000 0 0 $X=9272000 $Y=4968000
X2374 24 2348 dffr $T=9456000 9608000 1 180 $X=9272000 $Y=9608000
X2375 24 2349 dffr $T=9384000 1720000 0 0 $X=9384000 $Y=1720000
X2376 24 2350 dffr $T=9944000 10536000 1 180 $X=9760000 $Y=10536000
X2377 24 2351 dffr $T=10080000 8216000 1 180 $X=9896000 $Y=8216000
X2378 24 2352 dffr $T=10216000 5664000 1 180 $X=10032000 $Y=5664000
X2379 24 2353 dffr $T=10808000 3808000 1 180 $X=10624000 $Y=3808000
X2380 24 2268 dffr $T=10816000 328000 1 180 $X=10632000 $Y=328000
X2381 24 2354 dffr $T=10832000 560000 1 180 $X=10648000 $Y=560000
X2382 24 2355 dffr $T=11216000 8216000 0 0 $X=11216000 $Y=8216000
X2383 24 2356 dffr $T=11304000 3112000 0 0 $X=11304000 $Y=3112000
X2384 24 2357 dffr $T=11336000 8680000 0 0 $X=11336000 $Y=8680000
X2385 24 2358 dffr $T=12024000 9608000 1 180 $X=11840000 $Y=9608000
X2386 24 2359 dffr $T=11920000 7520000 0 0 $X=11920000 $Y=7520000
X2387 24 125 dffr $T=12192000 1720000 0 0 $X=12192000 $Y=1720000
X2388 24 2360 dffr $T=12264000 12624000 0 0 $X=12264000 $Y=12624000
X2389 24 178 dffr $T=12288000 1952000 0 0 $X=12288000 $Y=1952000
X2390 24 2361 dffr $T=12288000 11000000 0 0 $X=12288000 $Y=11000000
X2391 24 2362 dffr $T=12296000 3344000 0 0 $X=12296000 $Y=3344000
X2392 24 2363 dffr $T=12328000 10072000 0 0 $X=12328000 $Y=10072000
X2393 24 2364 dffr $T=12328000 11232000 0 0 $X=12328000 $Y=11232000
X2394 24 2365 dffr $T=12328000 12392000 0 0 $X=12328000 $Y=12392000
X2395 24 2366 dffr $T=12336000 5664000 0 0 $X=12336000 $Y=5664000
X2396 24 2367 dffr $T=12336000 13088000 0 0 $X=12336000 $Y=13088000
X2397 24 2368 dffr $T=12344000 2184000 0 0 $X=12344000 $Y=2184000
X2398 24 2369 dffr $T=12344000 2416000 0 0 $X=12344000 $Y=2416000
X2399 24 2370 dffr $T=12528000 2648000 1 180 $X=12344000 $Y=2648000
X2400 24 2371 dffr $T=12344000 3112000 0 0 $X=12344000 $Y=3112000
X2401 24 2372 dffr $T=12344000 3808000 0 0 $X=12344000 $Y=3808000
X2402 24 2373 dffr $T=12344000 4272000 0 0 $X=12344000 $Y=4272000
X2403 24 2374 dffr $T=12344000 4736000 0 0 $X=12344000 $Y=4736000
X2404 24 2375 dffr $T=12344000 4968000 0 0 $X=12344000 $Y=4968000
X2405 24 2376 dffr $T=12344000 5200000 0 0 $X=12344000 $Y=5200000
X2406 24 2377 dffr $T=12344000 5432000 0 0 $X=12344000 $Y=5432000
X2407 24 2378 dffr $T=12528000 6128000 1 180 $X=12344000 $Y=6128000
X2408 24 2379 dffr $T=12344000 6360000 0 0 $X=12344000 $Y=6360000
X2409 24 2380 dffr $T=12344000 6592000 0 0 $X=12344000 $Y=6592000
X2410 24 2381 dffr $T=12344000 7752000 0 0 $X=12344000 $Y=7752000
X2411 24 2382 dffr $T=12344000 7984000 0 0 $X=12344000 $Y=7984000
X2412 24 2383 dffr $T=12344000 8216000 0 0 $X=12344000 $Y=8216000
X2413 24 2384 dffr $T=12528000 8448000 1 180 $X=12344000 $Y=8448000
X2414 24 2385 dffr $T=12344000 9144000 0 0 $X=12344000 $Y=9144000
X2415 24 2386 dffr $T=12344000 9376000 0 0 $X=12344000 $Y=9376000
X2416 24 2387 dffr $T=12344000 9608000 0 0 $X=12344000 $Y=9608000
X2417 24 2388 dffr $T=12344000 9840000 0 0 $X=12344000 $Y=9840000
X2418 24 2389 dffr $T=12344000 10304000 0 0 $X=12344000 $Y=10304000
X2419 24 2390 dffr $T=12344000 10536000 0 0 $X=12344000 $Y=10536000
X2420 24 2391 dffr $T=12528000 10768000 1 180 $X=12344000 $Y=10768000
X2421 24 2392 dffr $T=12344000 11464000 0 0 $X=12344000 $Y=11464000
X2422 24 2393 dffr $T=12344000 11696000 0 0 $X=12344000 $Y=11696000
X2423 24 2394 dffr $T=12344000 11928000 0 0 $X=12344000 $Y=11928000
X2424 24 2395 dffr $T=12344000 12160000 0 0 $X=12344000 $Y=12160000
X2425 24 2396 dffr $T=12344000 12856000 0 0 $X=12344000 $Y=12856000
X2426 24 2397 inv01 $T=224000 3808000 0 0 $X=224000 $Y=3808000
X2427 24 2398 inv01 $T=344000 3576000 0 0 $X=344000 $Y=3576000
X2428 24 2399 inv01 $T=617000 3112000 1 180 $X=592000 $Y=3112000
X2429 24 2400 inv01 $T=728000 8912000 0 0 $X=728000 $Y=8912000
X2430 24 2401 inv01 $T=769000 3112000 1 180 $X=744000 $Y=3112000
X2431 24 2402 inv01 $T=785000 96000 1 180 $X=760000 $Y=96000
X2432 24 2403 inv01 $T=937000 2880000 1 180 $X=912000 $Y=2880000
X2433 24 2404 inv01 $T=1065000 560000 1 180 $X=1040000 $Y=560000
X2434 24 2405 inv01 $T=1233000 2648000 1 180 $X=1208000 $Y=2648000
X2435 24 2406 inv01 $T=1273000 1952000 1 180 $X=1248000 $Y=1952000
X2436 24 2407 inv01 $T=1393000 1256000 1 180 $X=1368000 $Y=1256000
X2437 24 2408 inv01 $T=1641000 1720000 1 180 $X=1616000 $Y=1720000
X2438 24 2409 inv01 $T=1673000 1720000 1 180 $X=1648000 $Y=1720000
X2439 24 2410 inv01 $T=1745000 1488000 1 180 $X=1720000 $Y=1488000
X2440 24 2411 inv01 $T=1745000 3112000 1 180 $X=1720000 $Y=3112000
X2441 24 2412 inv01 $T=1753000 2880000 1 180 $X=1728000 $Y=2880000
X2442 24 2413 inv01 $T=1769000 10072000 1 180 $X=1744000 $Y=10072000
X2443 24 2414 inv01 $T=1880000 10072000 0 0 $X=1880000 $Y=10072000
X2444 24 2415 inv01 $T=1944000 2416000 0 0 $X=1944000 $Y=2416000
X2445 24 2416 inv01 $T=2041000 2184000 1 180 $X=2016000 $Y=2184000
X2446 24 2417 inv01 $T=2128000 1488000 0 0 $X=2128000 $Y=1488000
X2447 24 2418 inv01 $T=2264000 3112000 0 0 $X=2264000 $Y=3112000
X2448 24 2419 inv01 $T=2377000 96000 1 180 $X=2352000 $Y=96000
X2449 24 2420 inv01 $T=2376000 3112000 0 0 $X=2376000 $Y=3112000
X2450 24 2421 inv01 $T=2529000 2648000 1 180 $X=2504000 $Y=2648000
X2451 24 2422 inv01 $T=2769000 2184000 1 180 $X=2744000 $Y=2184000
X2452 24 2423 inv01 $T=2777000 1488000 1 180 $X=2752000 $Y=1488000
X2453 24 2424 inv01 $T=2809000 2416000 1 180 $X=2784000 $Y=2416000
X2454 24 2425 inv01 $T=2841000 560000 1 180 $X=2816000 $Y=560000
X2455 24 2426 inv01 $T=2857000 96000 1 180 $X=2832000 $Y=96000
X2456 24 2427 inv01 $T=2993000 560000 1 180 $X=2968000 $Y=560000
X2457 24 2428 inv01 $T=2984000 328000 0 0 $X=2984000 $Y=328000
X2458 24 2429 inv01 $T=3049000 792000 1 180 $X=3024000 $Y=792000
X2459 24 2430 inv01 $T=3049000 1720000 1 180 $X=3024000 $Y=1720000
X2460 24 2431 inv01 $T=3065000 1256000 1 180 $X=3040000 $Y=1256000
X2461 24 2432 inv01 $T=3121000 96000 1 180 $X=3096000 $Y=96000
X2462 24 2433 inv01 $T=3153000 1488000 1 180 $X=3128000 $Y=1488000
X2463 24 2434 inv01 $T=3633000 96000 1 180 $X=3608000 $Y=96000
X2464 24 2435 inv01 $T=3616000 328000 0 0 $X=3616000 $Y=328000
X2465 24 2436 inv01 $T=3704000 96000 0 0 $X=3704000 $Y=96000
X2466 24 2437 inv01 $T=4072000 560000 0 0 $X=4072000 $Y=560000
X2467 24 2438 inv01 $T=4144000 96000 0 0 $X=4144000 $Y=96000
X2468 24 2439 inv01 $T=10729000 1488000 1 180 $X=10704000 $Y=1488000
X2469 24 2440 inv01 $T=10776000 1256000 0 0 $X=10776000 $Y=1256000
X2470 24 2354 inv01 $T=10832000 560000 0 0 $X=10832000 $Y=560000
X2471 24 2441 inv01 $T=10937000 328000 1 180 $X=10912000 $Y=328000
X2472 24 2442 inv01 $T=11192000 1488000 0 0 $X=11192000 $Y=1488000
X2473 24 2443 inv01 $T=11569000 1720000 1 180 $X=11544000 $Y=1720000
X2474 24 2444 inv01 $T=11657000 1488000 1 180 $X=11632000 $Y=1488000
X2475 24 2445 inv01 $T=11697000 6824000 1 180 $X=11672000 $Y=6824000
X2476 24 2446 inv01 $T=11793000 560000 1 180 $X=11768000 $Y=560000
X2477 24 2447 inv01 $T=11856000 7056000 0 0 $X=11856000 $Y=7056000
X2478 24 2448 inv01 $T=12096000 1720000 0 0 $X=12096000 $Y=1720000
X2479 24 2359 inv01 $T=12129000 7520000 1 180 $X=12104000 $Y=7520000
X2480 24 2449 inv01 $T=12273000 1488000 1 180 $X=12248000 $Y=1488000
X2481 24 2450 buf02 $T=185500 7752000 1 180 $X=152000 $Y=7752000
X2482 24 2451 buf02 $T=152000 9840000 0 0 $X=152000 $Y=9840000
X2483 24 2452 buf02 $T=152000 10072000 0 0 $X=152000 $Y=10072000
X2484 24 2453 buf02 $T=152000 12160000 0 0 $X=152000 $Y=12160000
X2485 24 2454 buf02 $T=225500 9840000 1 180 $X=192000 $Y=9840000
X2486 24 2455 buf02 $T=192000 10072000 0 0 $X=192000 $Y=10072000
X2487 24 2456 buf02 $T=192000 12160000 0 0 $X=192000 $Y=12160000
X2488 24 2457 buf02 $T=216000 11928000 0 0 $X=216000 $Y=11928000
X2489 24 2458 buf02 $T=400000 11464000 0 0 $X=400000 $Y=11464000
X2490 24 2459 buf02 $T=400000 12392000 0 0 $X=400000 $Y=12392000
X2491 24 2460 buf02 $T=400000 13320000 0 0 $X=400000 $Y=13320000
X2492 24 2461 buf02 $T=449500 9608000 1 180 $X=416000 $Y=9608000
X2493 24 2462 buf02 $T=456000 9608000 0 0 $X=456000 $Y=9608000
X2494 24 2463 buf02 $T=464000 7520000 0 0 $X=464000 $Y=7520000
X2495 24 2464 buf02 $T=464000 10304000 0 0 $X=464000 $Y=10304000
X2496 24 2465 buf02 $T=464000 13088000 0 0 $X=464000 $Y=13088000
X2497 24 2466 buf02 $T=504000 13320000 0 0 $X=504000 $Y=13320000
X2498 24 2467 buf02 $T=512000 10072000 0 0 $X=512000 $Y=10072000
X2499 24 2468 buf02 $T=512000 12160000 0 0 $X=512000 $Y=12160000
X2500 24 2469 buf02 $T=553500 9840000 1 180 $X=520000 $Y=9840000
X2501 24 2470 buf02 $T=553500 12624000 1 180 $X=520000 $Y=12624000
X2502 24 2471 buf02 $T=560000 9608000 0 0 $X=560000 $Y=9608000
X2503 24 2472 buf02 $T=593500 9840000 1 180 $X=560000 $Y=9840000
X2504 24 2289 buf02 $T=617500 9144000 1 180 $X=584000 $Y=9144000
X2505 24 2290 buf02 $T=617500 9376000 1 180 $X=584000 $Y=9376000
X2506 24 2473 buf02 $T=584000 10536000 0 0 $X=584000 $Y=10536000
X2507 24 2474 buf02 $T=584000 11696000 0 0 $X=584000 $Y=11696000
X2508 24 2475 buf02 $T=592000 10768000 0 0 $X=592000 $Y=10768000
X2509 24 2476 buf02 $T=633500 9840000 1 180 $X=600000 $Y=9840000
X2510 24 2477 buf02 $T=624000 9376000 0 0 $X=624000 $Y=9376000
X2511 24 2478 buf02 $T=632000 10768000 0 0 $X=632000 $Y=10768000
X2512 24 2479 buf02 $T=673500 9840000 1 180 $X=640000 $Y=9840000
X2513 24 2480 buf02 $T=648000 7984000 0 0 $X=648000 $Y=7984000
X2514 24 2481 buf02 $T=648000 12856000 0 0 $X=648000 $Y=12856000
X2515 24 2482 buf02 $T=697500 9376000 1 180 $X=664000 $Y=9376000
X2516 24 2483 buf02 $T=697500 11464000 1 180 $X=664000 $Y=11464000
X2517 24 2484 buf02 $T=705500 10072000 1 180 $X=672000 $Y=10072000
X2518 24 2485 buf02 $T=672000 11928000 0 0 $X=672000 $Y=11928000
X2519 24 2486 buf02 $T=680000 9840000 0 0 $X=680000 $Y=9840000
X2520 24 2487 buf02 $T=760000 7520000 0 0 $X=760000 $Y=7520000
X2521 24 2488 buf02 $T=801500 9376000 1 180 $X=768000 $Y=9376000
X2522 24 2489 buf02 $T=817500 7984000 1 180 $X=784000 $Y=7984000
X2523 24 2293 buf02 $T=784000 9608000 0 0 $X=784000 $Y=9608000
X2524 24 2490 buf02 $T=800000 7056000 0 0 $X=800000 $Y=7056000
X2525 24 2491 buf02 $T=833500 9144000 1 180 $X=800000 $Y=9144000
X2526 24 2492 buf02 $T=808000 9376000 0 0 $X=808000 $Y=9376000
X2527 24 2493 buf02 $T=816000 10304000 0 0 $X=816000 $Y=10304000
X2528 24 2494 buf02 $T=824000 11464000 0 0 $X=824000 $Y=11464000
X2529 24 2495 buf02 $T=857500 12160000 1 180 $X=824000 $Y=12160000
X2530 24 2496 buf02 $T=873500 9144000 1 180 $X=840000 $Y=9144000
X2531 24 2497 buf02 $T=864000 10072000 0 0 $X=864000 $Y=10072000
X2532 24 2498 buf02 $T=897500 12160000 1 180 $X=864000 $Y=12160000
X2533 24 2499 buf02 $T=921500 9608000 1 180 $X=888000 $Y=9608000
X2534 24 2500 buf02 $T=937500 12160000 1 180 $X=904000 $Y=12160000
X2535 24 2501 buf02 $T=945500 9144000 1 180 $X=912000 $Y=9144000
X2536 24 2502 buf02 $T=977500 9840000 1 180 $X=944000 $Y=9840000
X2537 24 2503 buf02 $T=993500 10072000 1 180 $X=960000 $Y=10072000
X2538 24 2504 buf02 $T=984000 9144000 0 0 $X=984000 $Y=9144000
X2539 24 2505 buf02 $T=1017500 9840000 1 180 $X=984000 $Y=9840000
X2540 24 2506 buf02 $T=984000 10768000 0 0 $X=984000 $Y=10768000
X2541 24 2507 buf02 $T=984000 11696000 0 0 $X=984000 $Y=11696000
X2542 24 2508 buf02 $T=992000 12624000 0 0 $X=992000 $Y=12624000
X2543 24 2509 buf02 $T=1000000 8680000 0 0 $X=1000000 $Y=8680000
X2544 24 2510 buf02 $T=1033500 12160000 1 180 $X=1000000 $Y=12160000
X2545 24 2511 buf02 $T=1024000 9144000 0 0 $X=1024000 $Y=9144000
X2546 24 2512 buf02 $T=1057500 9840000 1 180 $X=1024000 $Y=9840000
X2547 24 2513 buf02 $T=1057500 11696000 1 180 $X=1024000 $Y=11696000
X2548 24 2514 buf02 $T=1065500 12624000 1 180 $X=1032000 $Y=12624000
X2549 24 2515 buf02 $T=1089500 10072000 1 180 $X=1056000 $Y=10072000
X2550 24 2516 buf02 $T=1097500 9840000 1 180 $X=1064000 $Y=9840000
X2551 24 2517 buf02 $T=1105500 11928000 1 180 $X=1072000 $Y=11928000
X2552 24 2518 buf02 $T=1121500 12624000 1 180 $X=1088000 $Y=12624000
X2553 24 2519 buf02 $T=1129500 10072000 1 180 $X=1096000 $Y=10072000
X2554 24 2520 buf02 $T=1153500 9144000 1 180 $X=1120000 $Y=9144000
X2555 24 2521 buf02 $T=1120000 10536000 0 0 $X=1120000 $Y=10536000
X2556 24 2522 buf02 $T=1161500 9376000 1 180 $X=1128000 $Y=9376000
X2557 24 2523 buf02 $T=1193500 9144000 1 180 $X=1160000 $Y=9144000
X2558 24 2524 buf02 $T=1176000 12392000 0 0 $X=1176000 $Y=12392000
X2559 24 2525 buf02 $T=1257500 8448000 1 180 $X=1224000 $Y=8448000
X2560 24 2526 buf02 $T=1265500 9608000 1 180 $X=1232000 $Y=9608000
X2561 24 2527 buf02 $T=1256000 10072000 0 0 $X=1256000 $Y=10072000
X2562 24 2528 buf02 $T=1264000 11000000 0 0 $X=1264000 $Y=11000000
X2563 24 2529 buf02 $T=1305500 9608000 1 180 $X=1272000 $Y=9608000
X2564 24 2530 buf02 $T=1272000 12856000 0 0 $X=1272000 $Y=12856000
X2565 24 2531 buf02 $T=1321500 13320000 1 180 $X=1288000 $Y=13320000
X2566 24 2532 buf02 $T=1304000 11000000 0 0 $X=1304000 $Y=11000000
X2567 24 2533 buf02 $T=1345500 9608000 1 180 $X=1312000 $Y=9608000
X2568 24 2534 buf02 $T=1345500 12856000 1 180 $X=1312000 $Y=12856000
X2569 24 2535 buf02 $T=1328000 10072000 0 0 $X=1328000 $Y=10072000
X2570 24 2536 buf02 $T=1344000 11000000 0 0 $X=1344000 $Y=11000000
X2571 24 2537 buf02 $T=1385500 9608000 1 180 $X=1352000 $Y=9608000
X2572 24 2538 buf02 $T=1401500 10072000 1 180 $X=1368000 $Y=10072000
X2573 24 2539 buf02 $T=1384000 11000000 0 0 $X=1384000 $Y=11000000
X2574 24 2540 buf02 $T=1449500 7288000 1 180 $X=1416000 $Y=7288000
X2575 24 2541 buf02 $T=1448000 3112000 0 0 $X=1448000 $Y=3112000
X2576 24 2542 buf02 $T=1456000 13552000 0 0 $X=1456000 $Y=13552000
X2577 24 2543 buf02 $T=1521500 7288000 1 180 $X=1488000 $Y=7288000
X2578 24 2544 buf02 $T=1512000 8216000 0 0 $X=1512000 $Y=8216000
X2579 24 2545 buf02 $T=1545500 8448000 1 180 $X=1512000 $Y=8448000
X2580 24 2546 buf02 $T=1553500 7752000 1 180 $X=1520000 $Y=7752000
X2581 24 2547 buf02 $T=1528000 7288000 0 0 $X=1528000 $Y=7288000
X2582 24 2548 buf02 $T=1536000 12160000 0 0 $X=1536000 $Y=12160000
X2583 24 2549 buf02 $T=1585500 10536000 1 180 $X=1552000 $Y=10536000
X2584 24 2550 buf02 $T=1617500 8448000 1 180 $X=1584000 $Y=8448000
X2585 24 2551 buf02 $T=1633500 8912000 1 180 $X=1600000 $Y=8912000
X2586 24 2552 buf02 $T=1608000 8680000 0 0 $X=1608000 $Y=8680000
X2587 24 2553 buf02 $T=1608000 11696000 0 0 $X=1608000 $Y=11696000
X2588 24 2554 buf02 $T=1649500 9144000 1 180 $X=1616000 $Y=9144000
X2589 24 2555 buf02 $T=1665500 10304000 1 180 $X=1632000 $Y=10304000
X2590 24 2556 buf02 $T=1632000 12624000 0 0 $X=1632000 $Y=12624000
X2591 24 2557 buf02 $T=1681500 11696000 1 180 $X=1648000 $Y=11696000
X2592 24 2558 buf02 $T=1697500 10072000 1 180 $X=1664000 $Y=10072000
X2593 24 2559 buf02 $T=1713500 11928000 1 180 $X=1680000 $Y=11928000
X2594 24 2560 buf02 $T=1721500 11696000 1 180 $X=1688000 $Y=11696000
X2595 24 2561 buf02 $T=1745500 10536000 1 180 $X=1712000 $Y=10536000
X2596 24 2562 buf02 $T=1809500 11928000 1 180 $X=1776000 $Y=11928000
X2597 24 2563 buf02 $T=1817500 11696000 1 180 $X=1784000 $Y=11696000
X2598 24 2564 buf02 $T=1808000 2880000 0 0 $X=1808000 $Y=2880000
X2599 24 2565 buf02 $T=1816000 11928000 0 0 $X=1816000 $Y=11928000
X2600 24 2566 buf02 $T=1881500 2880000 1 180 $X=1848000 $Y=2880000
X2601 24 2567 buf02 $T=1848000 12856000 0 0 $X=1848000 $Y=12856000
X2602 24 2568 buf02 $T=1889500 11928000 1 180 $X=1856000 $Y=11928000
X2603 24 2569 buf02 $T=1936000 12392000 0 0 $X=1936000 $Y=12392000
X2604 24 2570 buf02 $T=2041500 11928000 1 180 $X=2008000 $Y=11928000
X2605 24 2571 buf02 $T=2048000 11000000 0 0 $X=2048000 $Y=11000000
X2606 24 2572 buf02 $T=2081500 11696000 1 180 $X=2048000 $Y=11696000
X2607 24 2573 buf02 $T=2089500 11232000 1 180 $X=2056000 $Y=11232000
X2608 24 2574 buf02 $T=2113500 12160000 1 180 $X=2080000 $Y=12160000
X2609 24 2575 buf02 $T=2121500 10072000 1 180 $X=2088000 $Y=10072000
X2610 24 2576 buf02 $T=2088000 11000000 0 0 $X=2088000 $Y=11000000
X2611 24 2577 buf02 $T=2096000 11232000 0 0 $X=2096000 $Y=11232000
X2612 24 2578 buf02 $T=2137500 10304000 1 180 $X=2104000 $Y=10304000
X2613 24 2579 buf02 $T=2120000 12160000 0 0 $X=2120000 $Y=12160000
X2614 24 2580 buf02 $T=2136000 12856000 0 0 $X=2136000 $Y=12856000
X2615 24 2581 buf02 $T=2160000 12160000 0 0 $X=2160000 $Y=12160000
X2616 24 2582 buf02 $T=2168000 10768000 0 0 $X=2168000 $Y=10768000
X2617 24 2583 buf02 $T=2225500 11000000 1 180 $X=2192000 $Y=11000000
X2618 24 2584 buf02 $T=2200000 12160000 0 0 $X=2200000 $Y=12160000
X2619 24 2585 buf02 $T=2280000 10536000 0 0 $X=2280000 $Y=10536000
X2620 24 2586 buf02 $T=2296000 11928000 0 0 $X=2296000 $Y=11928000
X2621 24 2587 buf02 $T=2345500 9144000 1 180 $X=2312000 $Y=9144000
X2622 24 2588 buf02 $T=2345500 13320000 1 180 $X=2312000 $Y=13320000
X2623 24 2589 buf02 $T=2353500 10304000 1 180 $X=2320000 $Y=10304000
X2624 24 2590 buf02 $T=2353500 10536000 1 180 $X=2320000 $Y=10536000
X2625 24 2591 buf02 $T=2344000 12392000 0 0 $X=2344000 $Y=12392000
X2626 24 2592 buf02 $T=2425500 10536000 1 180 $X=2392000 $Y=10536000
X2627 24 2593 buf02 $T=2449500 10304000 1 180 $X=2416000 $Y=10304000
X2628 24 2594 buf02 $T=2449500 11232000 1 180 $X=2416000 $Y=11232000
X2629 24 2595 buf02 $T=2457500 6824000 1 180 $X=2424000 $Y=6824000
X2630 24 2596 buf02 $T=2440000 12856000 0 0 $X=2440000 $Y=12856000
X2631 24 2597 buf02 $T=2481500 8680000 1 180 $X=2448000 $Y=8680000
X2632 24 2598 buf02 $T=2489500 10768000 1 180 $X=2456000 $Y=10768000
X2633 24 2599 buf02 $T=2488000 12160000 0 0 $X=2488000 $Y=12160000
X2634 24 2600 buf02 $T=2537500 1720000 1 180 $X=2504000 $Y=1720000
X2635 24 2601 buf02 $T=2561500 12160000 1 180 $X=2528000 $Y=12160000
X2636 24 2602 buf02 $T=2577500 11928000 1 180 $X=2544000 $Y=11928000
X2637 24 2603 buf02 $T=2568000 12160000 0 0 $X=2568000 $Y=12160000
X2638 24 2604 buf02 $T=2641500 12160000 1 180 $X=2608000 $Y=12160000
X2639 24 2605 buf02 $T=2608000 12856000 0 0 $X=2608000 $Y=12856000
X2640 24 2606 buf02 $T=2657500 10304000 1 180 $X=2624000 $Y=10304000
X2641 24 2607 buf02 $T=2697500 10304000 1 180 $X=2664000 $Y=10304000
X2642 24 2608 buf02 $T=2705500 9376000 1 180 $X=2672000 $Y=9376000
X2643 24 2609 buf02 $T=2696000 12392000 0 0 $X=2696000 $Y=12392000
X2644 24 2610 buf02 $T=2729500 12624000 1 180 $X=2696000 $Y=12624000
X2645 24 2611 buf02 $T=2712000 6824000 0 0 $X=2712000 $Y=6824000
X2646 24 2612 buf02 $T=2769500 11464000 1 180 $X=2736000 $Y=11464000
X2647 24 2613 buf02 $T=2793500 11928000 1 180 $X=2760000 $Y=11928000
X2648 24 2614 buf02 $T=2801500 1952000 1 180 $X=2768000 $Y=1952000
X2649 24 2615 buf02 $T=2776000 11464000 0 0 $X=2776000 $Y=11464000
X2650 24 2616 buf02 $T=2809500 11696000 1 180 $X=2776000 $Y=11696000
X2651 24 2617 buf02 $T=2784000 11000000 0 0 $X=2784000 $Y=11000000
X2652 24 2618 buf02 $T=2832000 13320000 0 0 $X=2832000 $Y=13320000
X2653 24 2619 buf02 $T=2832000 13552000 0 0 $X=2832000 $Y=13552000
X2654 24 2620 buf02 $T=2881500 7288000 1 180 $X=2848000 $Y=7288000
X2655 24 2621 buf02 $T=2897500 10768000 1 180 $X=2864000 $Y=10768000
X2656 24 2622 buf02 $T=2880000 2416000 0 0 $X=2880000 $Y=2416000
X2657 24 2623 buf02 $T=2921500 13088000 1 180 $X=2888000 $Y=13088000
X2658 24 2624 buf02 $T=2937500 11464000 1 180 $X=2904000 $Y=11464000
X2659 24 2625 buf02 $T=2928000 11696000 0 0 $X=2928000 $Y=11696000
X2660 24 2626 buf02 $T=2936000 11232000 0 0 $X=2936000 $Y=11232000
X2661 24 2627 buf02 $T=2977500 11464000 1 180 $X=2944000 $Y=11464000
X2662 24 2628 buf02 $T=2968000 12856000 0 0 $X=2968000 $Y=12856000
X2663 24 2629 buf02 $T=3009500 11232000 1 180 $X=2976000 $Y=11232000
X2664 24 2630 buf02 $T=2984000 12392000 0 0 $X=2984000 $Y=12392000
X2665 24 2631 buf02 $T=3016000 11232000 0 0 $X=3016000 $Y=11232000
X2666 24 2632 buf02 $T=3048000 9376000 0 0 $X=3048000 $Y=9376000
X2667 24 2633 buf02 $T=3089500 11000000 1 180 $X=3056000 $Y=11000000
X2668 24 2634 buf02 $T=3089500 11232000 1 180 $X=3056000 $Y=11232000
X2669 24 2635 buf02 $T=3080000 11696000 0 0 $X=3080000 $Y=11696000
X2670 24 2636 buf02 $T=3129500 11232000 1 180 $X=3096000 $Y=11232000
X2671 24 2637 buf02 $T=3137500 10072000 1 180 $X=3104000 $Y=10072000
X2672 24 2638 buf02 $T=3153500 11696000 1 180 $X=3120000 $Y=11696000
X2673 24 2639 buf02 $T=3169500 11232000 1 180 $X=3136000 $Y=11232000
X2674 24 2640 buf02 $T=3193500 11696000 1 180 $X=3160000 $Y=11696000
X2675 24 2641 buf02 $T=3217500 12160000 1 180 $X=3184000 $Y=12160000
X2676 24 2642 buf02 $T=3225500 10768000 1 180 $X=3192000 $Y=10768000
X2677 24 2643 buf02 $T=3233500 11696000 1 180 $X=3200000 $Y=11696000
X2678 24 2644 buf02 $T=3257500 12160000 1 180 $X=3224000 $Y=12160000
X2679 24 2645 buf02 $T=3432000 12160000 0 0 $X=3432000 $Y=12160000
X2680 24 2646 buf02 $T=3472000 12160000 0 0 $X=3472000 $Y=12160000
X2681 24 2647 buf02 $T=3488000 9144000 0 0 $X=3488000 $Y=9144000
X2682 24 2648 buf02 $T=3545500 10072000 1 180 $X=3512000 $Y=10072000
X2683 24 2649 buf02 $T=3640000 9376000 0 0 $X=3640000 $Y=9376000
X2684 24 2650 buf02 $T=3697500 10072000 1 180 $X=3664000 $Y=10072000
X2685 24 2651 buf02 $T=3672000 13088000 0 0 $X=3672000 $Y=13088000
X2686 24 2652 buf02 $T=3680000 13552000 0 0 $X=3680000 $Y=13552000
X2687 24 2653 buf02 $T=3704000 10072000 0 0 $X=3704000 $Y=10072000
X2688 24 2654 buf02 $T=3720000 13552000 0 0 $X=3720000 $Y=13552000
X2689 24 2655 buf02 $T=3752000 13320000 0 0 $X=3752000 $Y=13320000
X2690 24 2656 buf02 $T=3760000 12624000 0 0 $X=3760000 $Y=12624000
X2691 24 2657 buf02 $T=3768000 13088000 0 0 $X=3768000 $Y=13088000
X2692 24 2658 buf02 $T=3809500 11928000 1 180 $X=3776000 $Y=11928000
X2693 24 2659 buf02 $T=3905500 9840000 1 180 $X=3872000 $Y=9840000
X2694 24 2660 buf02 $T=3937500 10304000 1 180 $X=3904000 $Y=10304000
X2695 24 2661 buf02 $T=3945500 9840000 1 180 $X=3912000 $Y=9840000
X2696 24 2662 buf02 $T=3985500 10536000 1 180 $X=3952000 $Y=10536000
X2697 24 2663 buf02 $T=4025500 9144000 1 180 $X=3992000 $Y=9144000
X2698 24 2664 buf02 $T=3992000 10072000 0 0 $X=3992000 $Y=10072000
X2699 24 2665 buf02 $T=4008000 13552000 0 0 $X=4008000 $Y=13552000
X2700 24 2666 buf02 $T=4024000 12160000 0 0 $X=4024000 $Y=12160000
X2701 24 2667 buf02 $T=4032000 9144000 0 0 $X=4032000 $Y=9144000
X2702 24 2668 buf02 $T=4048000 10768000 0 0 $X=4048000 $Y=10768000
X2703 24 2669 buf02 $T=4081500 12856000 1 180 $X=4048000 $Y=12856000
X2704 24 2670 buf02 $T=4081500 13552000 1 180 $X=4048000 $Y=13552000
X2705 24 2671 buf02 $T=4096000 13320000 0 0 $X=4096000 $Y=13320000
X2706 24 2672 buf02 $T=4177500 13552000 1 180 $X=4144000 $Y=13552000
X2707 24 2673 buf02 $T=4193500 12624000 1 180 $X=4160000 $Y=12624000
X2708 24 2674 buf02 $T=4225500 13320000 1 180 $X=4192000 $Y=13320000
X2709 24 2675 buf02 $T=4265500 12624000 1 180 $X=4232000 $Y=12624000
X2710 24 2676 buf02 $T=4273500 13552000 1 180 $X=4240000 $Y=13552000
X2711 24 2677 buf02 $T=4256000 11464000 0 0 $X=4256000 $Y=11464000
X2712 24 2678 buf02 $T=4376000 11232000 0 0 $X=4376000 $Y=11232000
X2713 24 2679 buf02 $T=4392000 12392000 0 0 $X=4392000 $Y=12392000
X2714 24 2680 buf02 $T=4433500 11928000 1 180 $X=4400000 $Y=11928000
X2715 24 2681 buf02 $T=4424000 10536000 0 0 $X=4424000 $Y=10536000
X2716 24 2682 buf02 $T=4465500 9144000 1 180 $X=4432000 $Y=9144000
X2717 24 2683 buf02 $T=4465500 12392000 1 180 $X=4432000 $Y=12392000
X2718 24 2684 buf02 $T=4504000 12160000 0 0 $X=4504000 $Y=12160000
X2719 24 2685 buf02 $T=4528000 10536000 0 0 $X=4528000 $Y=10536000
X2720 24 2686 buf02 $T=4536000 10768000 0 0 $X=4536000 $Y=10768000
X2721 24 2687 buf02 $T=4577500 12160000 1 180 $X=4544000 $Y=12160000
X2722 24 2688 buf02 $T=4593500 10072000 1 180 $X=4560000 $Y=10072000
X2723 24 2689 buf02 $T=4600000 11464000 0 0 $X=4600000 $Y=11464000
X2724 24 2690 buf02 $T=4649500 12160000 1 180 $X=4616000 $Y=12160000
X2725 24 2691 buf02 $T=4657500 10304000 1 180 $X=4624000 $Y=10304000
X2726 24 2692 buf02 $T=4689500 12160000 1 180 $X=4656000 $Y=12160000
X2727 24 2693 buf02 $T=4729500 7752000 1 180 $X=4696000 $Y=7752000
X2728 24 2694 buf02 $T=4729500 8216000 1 180 $X=4696000 $Y=8216000
X2729 24 2695 buf02 $T=4720000 11232000 0 0 $X=4720000 $Y=11232000
X2730 24 2696 buf02 $T=4769500 8216000 1 180 $X=4736000 $Y=8216000
X2731 24 2697 buf02 $T=4760000 11232000 0 0 $X=4760000 $Y=11232000
X2732 24 2698 buf02 $T=4784000 11696000 0 0 $X=4784000 $Y=11696000
X2733 24 2699 buf02 $T=4881500 13088000 1 180 $X=4848000 $Y=13088000
X2734 24 2700 buf02 $T=4913500 10072000 1 180 $X=4880000 $Y=10072000
X2735 24 2701 buf02 $T=4920000 12392000 0 0 $X=4920000 $Y=12392000
X2736 24 2702 buf02 $T=4977500 13088000 1 180 $X=4944000 $Y=13088000
X2737 24 2703 buf02 $T=4960000 13552000 0 0 $X=4960000 $Y=13552000
X2738 24 2704 buf02 $T=5064000 13552000 0 0 $X=5064000 $Y=13552000
X2739 24 2705 buf02 $T=5080000 10536000 0 0 $X=5080000 $Y=10536000
X2740 24 2706 buf02 $T=5080000 12392000 0 0 $X=5080000 $Y=12392000
X2741 24 2707 buf02 $T=5080000 12624000 0 0 $X=5080000 $Y=12624000
X2742 24 2708 buf02 $T=5104000 11232000 0 0 $X=5104000 $Y=11232000
X2743 24 2709 buf02 $T=5104000 11696000 0 0 $X=5104000 $Y=11696000
X2744 24 2710 buf02 $T=5112000 11000000 0 0 $X=5112000 $Y=11000000
X2745 24 2711 buf02 $T=5153500 12856000 1 180 $X=5120000 $Y=12856000
X2746 24 2712 buf02 $T=5144000 11232000 0 0 $X=5144000 $Y=11232000
X2747 24 2713 buf02 $T=5144000 11696000 0 0 $X=5144000 $Y=11696000
X2748 24 2714 buf02 $T=5201500 10072000 1 180 $X=5168000 $Y=10072000
X2749 24 2715 buf02 $T=5209500 12392000 1 180 $X=5176000 $Y=12392000
X2750 24 2716 buf02 $T=5241500 10072000 1 180 $X=5208000 $Y=10072000
X2751 24 2717 buf02 $T=5208000 10536000 0 0 $X=5208000 $Y=10536000
X2752 24 2718 buf02 $T=5273500 10304000 1 180 $X=5240000 $Y=10304000
X2753 24 2719 buf02 $T=5240000 11000000 0 0 $X=5240000 $Y=11000000
X2754 24 2720 buf02 $T=5281500 11464000 1 180 $X=5248000 $Y=11464000
X2755 24 2721 buf02 $T=5281500 12392000 1 180 $X=5248000 $Y=12392000
X2756 24 2722 buf02 $T=5289500 12160000 1 180 $X=5256000 $Y=12160000
X2757 24 2723 buf02 $T=5321500 11232000 1 180 $X=5288000 $Y=11232000
X2758 24 2724 buf02 $T=5329500 11928000 1 180 $X=5296000 $Y=11928000
X2759 24 2725 buf02 $T=5329500 12160000 1 180 $X=5296000 $Y=12160000
X2760 24 2726 buf02 $T=5337500 10536000 1 180 $X=5304000 $Y=10536000
X2761 24 2727 buf02 $T=5345500 9376000 1 180 $X=5312000 $Y=9376000
X2762 24 2728 buf02 $T=5401500 11000000 1 180 $X=5368000 $Y=11000000
X2763 24 2729 buf02 $T=5417500 12624000 1 180 $X=5384000 $Y=12624000
X2764 24 2730 buf02 $T=5425500 9608000 1 180 $X=5392000 $Y=9608000
X2765 24 2731 buf02 $T=5392000 10304000 0 0 $X=5392000 $Y=10304000
X2766 24 2732 buf02 $T=5465500 10304000 1 180 $X=5432000 $Y=10304000
X2767 24 2733 buf02 $T=5545500 13320000 1 180 $X=5512000 $Y=13320000
X2768 24 2734 buf02 $T=5577500 13088000 1 180 $X=5544000 $Y=13088000
X2769 24 2735 buf02 $T=5552000 11696000 0 0 $X=5552000 $Y=11696000
X2770 24 2736 buf02 $T=5560000 10072000 0 0 $X=5560000 $Y=10072000
X2771 24 2737 buf02 $T=5593500 10304000 1 180 $X=5560000 $Y=10304000
X2772 24 2324 buf02 $T=5609500 11928000 1 180 $X=5576000 $Y=11928000
X2773 24 2738 buf02 $T=5633500 9376000 1 180 $X=5600000 $Y=9376000
X2774 24 2739 buf02 $T=5600000 10768000 0 0 $X=5600000 $Y=10768000
X2775 24 2740 buf02 $T=5673500 9376000 1 180 $X=5640000 $Y=9376000
X2776 24 2741 buf02 $T=5697500 8448000 1 180 $X=5664000 $Y=8448000
X2777 24 2742 buf02 $T=5672000 11232000 0 0 $X=5672000 $Y=11232000
X2778 24 2743 buf02 $T=5737500 12392000 1 180 $X=5704000 $Y=12392000
X2779 24 2744 buf02 $T=5712000 11232000 0 0 $X=5712000 $Y=11232000
X2780 24 2745 buf02 $T=5720000 13552000 0 0 $X=5720000 $Y=13552000
X2781 24 2746 buf02 $T=5769500 9608000 1 180 $X=5736000 $Y=9608000
X2782 24 2747 buf02 $T=5793500 12624000 1 180 $X=5760000 $Y=12624000
X2783 24 2748 buf02 $T=5801500 8448000 1 180 $X=5768000 $Y=8448000
X2784 24 2749 buf02 $T=5768000 10536000 0 0 $X=5768000 $Y=10536000
X2785 24 2750 buf02 $T=5808000 11232000 0 0 $X=5808000 $Y=11232000
X2786 24 2751 buf02 $T=5840000 11464000 0 0 $X=5840000 $Y=11464000
X2787 24 2752 buf02 $T=5897500 13088000 1 180 $X=5864000 $Y=13088000
X2788 24 2753 buf02 $T=5905500 13320000 1 180 $X=5872000 $Y=13320000
X2789 24 2754 buf02 $T=6000000 11232000 0 0 $X=6000000 $Y=11232000
X2790 24 2755 buf02 $T=6065500 10072000 1 180 $X=6032000 $Y=10072000
X2791 24 2756 buf02 $T=6065500 13320000 1 180 $X=6032000 $Y=13320000
X2792 24 2757 buf02 $T=6073500 11232000 1 180 $X=6040000 $Y=11232000
X2793 24 2758 buf02 $T=6073500 11696000 1 180 $X=6040000 $Y=11696000
X2794 24 2759 buf02 $T=6081500 10768000 1 180 $X=6048000 $Y=10768000
X2795 24 2760 buf02 $T=6081500 11928000 1 180 $X=6048000 $Y=11928000
X2796 24 2761 buf02 $T=6097500 11464000 1 180 $X=6064000 $Y=11464000
X2797 24 2762 buf02 $T=6105500 10072000 1 180 $X=6072000 $Y=10072000
X2798 24 2763 buf02 $T=6121500 10768000 1 180 $X=6088000 $Y=10768000
X2799 24 2764 buf02 $T=6121500 12392000 1 180 $X=6088000 $Y=12392000
X2800 24 2765 buf02 $T=6104000 10304000 0 0 $X=6104000 $Y=10304000
X2801 24 2766 buf02 $T=6153500 10536000 1 180 $X=6120000 $Y=10536000
X2802 24 2767 buf02 $T=6177500 10304000 1 180 $X=6144000 $Y=10304000
X2803 24 2768 buf02 $T=6185500 8448000 1 180 $X=6152000 $Y=8448000
X2804 24 2769 buf02 $T=6185500 9376000 1 180 $X=6152000 $Y=9376000
X2805 24 2770 buf02 $T=6225500 8448000 1 180 $X=6192000 $Y=8448000
X2806 24 2771 buf02 $T=6241500 9840000 1 180 $X=6208000 $Y=9840000
X2807 24 2772 buf02 $T=6297500 8448000 1 180 $X=6264000 $Y=8448000
X2808 24 2773 buf02 $T=6313500 9840000 1 180 $X=6280000 $Y=9840000
X2809 24 2328 buf02 $T=6296000 10072000 0 0 $X=6296000 $Y=10072000
X2810 24 2774 buf02 $T=6369500 10072000 1 180 $X=6336000 $Y=10072000
X2811 24 2775 buf02 $T=6400000 13088000 0 0 $X=6400000 $Y=13088000
X2812 24 2776 buf02 $T=6441500 10072000 1 180 $X=6408000 $Y=10072000
X2813 24 2777 buf02 $T=7337500 9144000 1 180 $X=7304000 $Y=9144000
X2814 24 2778 buf02 $T=7304000 11232000 0 0 $X=7304000 $Y=11232000
X2815 24 2779 buf02 $T=7337500 11464000 1 180 $X=7304000 $Y=11464000
X2816 24 2780 buf02 $T=7337500 11696000 1 180 $X=7304000 $Y=11696000
X2817 24 2781 buf02 $T=7441500 11232000 1 180 $X=7408000 $Y=11232000
X2818 24 2782 buf02 $T=7784000 11928000 0 0 $X=7784000 $Y=11928000
X2819 24 2783 buf02 $T=7841500 11696000 1 180 $X=7808000 $Y=11696000
X2820 24 2784 buf02 $T=7872000 9840000 0 0 $X=7872000 $Y=9840000
X2821 24 2785 buf02 $T=7896000 11464000 0 0 $X=7896000 $Y=11464000
X2822 24 2786 buf02 $T=7936000 9608000 0 0 $X=7936000 $Y=9608000
X2823 24 2787 buf02 $T=7944000 11232000 0 0 $X=7944000 $Y=11232000
X2824 24 2788 buf02 $T=8056000 13088000 0 0 $X=8056000 $Y=13088000
X2825 24 2789 buf02 $T=8088000 13552000 0 0 $X=8088000 $Y=13552000
X2826 24 2790 buf02 $T=8160000 13088000 0 0 $X=8160000 $Y=13088000
X2827 24 2791 buf02 $T=8264000 13320000 0 0 $X=8264000 $Y=13320000
X2828 24 2792 buf02 $T=8480000 13088000 0 0 $X=8480000 $Y=13088000
X2829 24 2793 buf02 $T=8569500 11928000 1 180 $X=8536000 $Y=11928000
X2830 24 2794 buf02 $T=8568000 12856000 0 0 $X=8568000 $Y=12856000
X2831 24 2795 buf02 $T=8792000 11696000 0 0 $X=8792000 $Y=11696000
X2832 24 2796 buf02 $T=8832000 12160000 0 0 $X=8832000 $Y=12160000
X2833 24 2797 buf02 $T=8872000 11928000 0 0 $X=8872000 $Y=11928000
X2834 24 2798 buf02 $T=8945500 10072000 1 180 $X=8912000 $Y=10072000
X2835 24 2799 buf02 $T=8952000 10072000 0 0 $X=8952000 $Y=10072000
X2836 24 2800 buf02 $T=9009500 11464000 1 180 $X=8976000 $Y=11464000
X2837 24 2801 buf02 $T=8984000 12624000 0 0 $X=8984000 $Y=12624000
X2838 24 2802 buf02 $T=9056000 10072000 0 0 $X=9056000 $Y=10072000
X2839 24 2803 buf02 $T=9056000 12624000 0 0 $X=9056000 $Y=12624000
X2840 24 2804 buf02 $T=9105500 11928000 1 180 $X=9072000 $Y=11928000
X2841 24 2805 buf02 $T=9096000 10072000 0 0 $X=9096000 $Y=10072000
X2842 24 2806 buf02 $T=9096000 11232000 0 0 $X=9096000 $Y=11232000
X2843 24 2807 buf02 $T=9136000 10072000 0 0 $X=9136000 $Y=10072000
X2844 24 2808 buf02 $T=9136000 11464000 0 0 $X=9136000 $Y=11464000
X2845 24 2809 buf02 $T=9176000 10072000 0 0 $X=9176000 $Y=10072000
X2846 24 2810 buf02 $T=9225500 11232000 1 180 $X=9192000 $Y=11232000
X2847 24 2811 buf02 $T=9216000 10072000 0 0 $X=9216000 $Y=10072000
X2848 24 2812 buf02 $T=9265500 11464000 1 180 $X=9232000 $Y=11464000
X2849 24 2813 buf02 $T=9344000 12624000 0 0 $X=9344000 $Y=12624000
X2850 24 2814 buf02 $T=9368000 13552000 0 0 $X=9368000 $Y=13552000
X2851 24 2815 buf02 $T=9376000 13088000 0 0 $X=9376000 $Y=13088000
X2852 24 2816 buf02 $T=9417500 12624000 1 180 $X=9384000 $Y=12624000
X2853 24 2817 buf02 $T=9400000 12856000 0 0 $X=9400000 $Y=12856000
X2854 24 2818 buf02 $T=9408000 13552000 0 0 $X=9408000 $Y=13552000
X2855 24 2819 buf02 $T=9416000 13088000 0 0 $X=9416000 $Y=13088000
X2856 24 2820 buf02 $T=9489500 13088000 1 180 $X=9456000 $Y=13088000
X2857 24 2821 buf02 $T=9480000 12392000 0 0 $X=9480000 $Y=12392000
X2858 24 2822 buf02 $T=9488000 12160000 0 0 $X=9488000 $Y=12160000
X2859 24 2823 buf02 $T=9496000 12856000 0 0 $X=9496000 $Y=12856000
X2860 24 2824 buf02 $T=9553500 12392000 1 180 $X=9520000 $Y=12392000
X2861 24 2825 buf02 $T=9569500 12856000 1 180 $X=9536000 $Y=12856000
X2862 24 2826 buf02 $T=9617500 13088000 1 180 $X=9584000 $Y=13088000
X2863 24 2827 buf02 $T=9592000 12392000 0 0 $X=9592000 $Y=12392000
X2864 24 2828 buf02 $T=9665500 12392000 1 180 $X=9632000 $Y=12392000
X2865 24 2829 buf02 $T=9705500 12392000 1 180 $X=9672000 $Y=12392000
X2866 24 2830 buf02 $T=9680000 9144000 0 0 $X=9680000 $Y=9144000
X2867 24 2831 buf02 $T=9713500 13088000 1 180 $X=9680000 $Y=13088000
X2868 24 2832 buf02 $T=9721500 12856000 1 180 $X=9688000 $Y=12856000
X2869 24 2833 buf02 $T=9696000 11928000 0 0 $X=9696000 $Y=11928000
X2870 24 2834 buf02 $T=9753500 13088000 1 180 $X=9720000 $Y=13088000
X2871 24 2835 buf02 $T=9761500 12856000 1 180 $X=9728000 $Y=12856000
X2872 24 2836 buf02 $T=9728000 13552000 0 0 $X=9728000 $Y=13552000
X2873 24 2837 buf02 $T=9760000 13320000 0 0 $X=9760000 $Y=13320000
X2874 24 2838 buf02 $T=9768000 13552000 0 0 $X=9768000 $Y=13552000
X2875 24 2839 buf02 $T=9792000 11464000 0 0 $X=9792000 $Y=11464000
X2876 24 2840 buf02 $T=9800000 13320000 0 0 $X=9800000 $Y=13320000
X2877 24 2841 buf02 $T=9841500 13552000 1 180 $X=9808000 $Y=13552000
X2878 24 2842 buf02 $T=9816000 12624000 0 0 $X=9816000 $Y=12624000
X2879 24 2843 buf02 $T=9873500 8912000 1 180 $X=9840000 $Y=8912000
X2880 24 2844 buf02 $T=9881500 11928000 1 180 $X=9848000 $Y=11928000
X2881 24 2845 buf02 $T=9856000 11696000 0 0 $X=9856000 $Y=11696000
X2882 24 2846 buf02 $T=9856000 12624000 0 0 $X=9856000 $Y=12624000
X2883 24 2847 buf02 $T=9872000 12160000 0 0 $X=9872000 $Y=12160000
X2884 24 2848 buf02 $T=9880000 8912000 0 0 $X=9880000 $Y=8912000
X2885 24 2849 buf02 $T=9961500 13088000 1 180 $X=9928000 $Y=13088000
X2886 24 2850 buf02 $T=10017500 12624000 1 180 $X=9984000 $Y=12624000
X2887 24 2851 buf02 $T=10000000 12856000 0 0 $X=10000000 $Y=12856000
X2888 24 2852 buf02 $T=10032000 12160000 0 0 $X=10032000 $Y=12160000
X2889 24 2853 buf02 $T=10105500 12160000 1 180 $X=10072000 $Y=12160000
X2890 24 2854 buf02 $T=10144000 13320000 0 0 $X=10144000 $Y=13320000
X2891 24 2855 buf02 $T=10201500 13088000 1 180 $X=10168000 $Y=13088000
X2892 24 2856 buf02 $T=10184000 13320000 0 0 $X=10184000 $Y=13320000
X2893 24 2857 buf02 $T=10224000 13320000 0 0 $X=10224000 $Y=13320000
X2894 24 2858 buf02 $T=10296000 11696000 0 0 $X=10296000 $Y=11696000
X2895 24 2859 buf02 $T=10329500 13088000 1 180 $X=10296000 $Y=13088000
X2896 24 2860 buf02 $T=10361500 12856000 1 180 $X=10328000 $Y=12856000
X2897 24 2861 buf02 $T=10369500 12624000 1 180 $X=10336000 $Y=12624000
X2898 24 2862 buf02 $T=10369500 13088000 1 180 $X=10336000 $Y=13088000
X2899 24 2863 buf02 $T=10344000 9608000 0 0 $X=10344000 $Y=9608000
X2900 24 2864 buf02 $T=10368000 12856000 0 0 $X=10368000 $Y=12856000
X2901 24 2865 buf02 $T=10409500 12624000 1 180 $X=10376000 $Y=12624000
X2902 24 2866 buf02 $T=10384000 11464000 0 0 $X=10384000 $Y=11464000
X2903 24 2867 buf02 $T=10425500 10072000 1 180 $X=10392000 $Y=10072000
X2904 24 2868 buf02 $T=10408000 12856000 0 0 $X=10408000 $Y=12856000
X2905 24 2869 buf02 $T=10449500 12624000 1 180 $X=10416000 $Y=12624000
X2906 24 2870 buf02 $T=10440000 13088000 0 0 $X=10440000 $Y=13088000
X2907 24 2871 buf02 $T=10481500 12856000 1 180 $X=10448000 $Y=12856000
X2908 24 2872 buf02 $T=10489500 12624000 1 180 $X=10456000 $Y=12624000
X2909 24 2873 buf02 $T=10496000 12624000 0 0 $X=10496000 $Y=12624000
X2910 24 2874 buf02 $T=10600000 11464000 0 0 $X=10600000 $Y=11464000
X2911 24 2875 buf02 $T=10633500 12624000 1 180 $X=10600000 $Y=12624000
X2912 24 2876 buf02 $T=10760000 3112000 0 0 $X=10760000 $Y=3112000
X2913 24 2877 buf02 $T=10840000 10072000 0 0 $X=10840000 $Y=10072000
X2914 24 2878 buf02 $T=10888000 11464000 0 0 $X=10888000 $Y=11464000
X2915 24 2879 buf02 $T=10952000 13088000 0 0 $X=10952000 $Y=13088000
X2916 24 2880 buf02 $T=11081500 12160000 1 180 $X=11048000 $Y=12160000
X2917 24 2881 buf02 $T=11048000 13088000 0 0 $X=11048000 $Y=13088000
X2918 24 2882 buf02 $T=11137500 12624000 1 180 $X=11104000 $Y=12624000
X2919 24 2883 buf02 $T=11145500 12392000 1 180 $X=11112000 $Y=12392000
X2920 24 2884 buf02 $T=11177500 12624000 1 180 $X=11144000 $Y=12624000
X2921 24 2885 buf02 $T=11185500 13088000 1 180 $X=11152000 $Y=13088000
X2922 24 2886 buf02 $T=11201500 10072000 1 180 $X=11168000 $Y=10072000
X2923 24 2887 buf02 $T=11225500 13088000 1 180 $X=11192000 $Y=13088000
X2924 24 2888 buf02 $T=11273500 12624000 1 180 $X=11240000 $Y=12624000
X2925 24 2889 buf02 $T=11256000 13552000 0 0 $X=11256000 $Y=13552000
X2926 24 2890 buf02 $T=11280000 12624000 0 0 $X=11280000 $Y=12624000
X2927 24 2891 buf02 $T=11353500 12624000 1 180 $X=11320000 $Y=12624000
X2928 24 2892 buf02 $T=11376000 9608000 0 0 $X=11376000 $Y=9608000
X2929 24 2893 buf02 $T=11425500 12624000 1 180 $X=11392000 $Y=12624000
X2930 24 2894 buf02 $T=11433500 1488000 1 180 $X=11400000 $Y=1488000
X2931 24 2895 buf02 $T=11441500 12160000 1 180 $X=11408000 $Y=12160000
X2932 24 2896 buf02 $T=11465500 13320000 1 180 $X=11432000 $Y=13320000
X2933 24 2897 buf02 $T=11473500 1488000 1 180 $X=11440000 $Y=1488000
X2934 24 2898 buf02 $T=11489500 10072000 1 180 $X=11456000 $Y=10072000
X2935 24 2899 buf02 $T=11504000 13320000 0 0 $X=11504000 $Y=13320000
X2936 24 2900 buf02 $T=11544000 13320000 0 0 $X=11544000 $Y=13320000
X2937 24 2901 buf02 $T=11585500 12856000 1 180 $X=11552000 $Y=12856000
X2938 24 2902 buf02 $T=11617500 13320000 1 180 $X=11584000 $Y=13320000
X2939 24 2903 buf02 $T=11600000 13088000 0 0 $X=11600000 $Y=13088000
X2940 24 2904 buf02 $T=11657500 13320000 1 180 $X=11624000 $Y=13320000
X2941 24 2905 buf02 $T=11648000 12856000 0 0 $X=11648000 $Y=12856000
X2942 24 2906 buf02 $T=11697500 13320000 1 180 $X=11664000 $Y=13320000
X2943 24 2907 buf02 $T=11688000 12160000 0 0 $X=11688000 $Y=12160000
X2944 24 2908 buf02 $T=11721500 12392000 1 180 $X=11688000 $Y=12392000
X2945 24 2909 buf02 $T=11688000 12856000 0 0 $X=11688000 $Y=12856000
X2946 24 2910 buf02 $T=11793500 12856000 1 180 $X=11760000 $Y=12856000
X2947 24 2911 buf02 $T=11832000 12624000 0 0 $X=11832000 $Y=12624000
X2948 24 2912 buf02 $T=11872000 12624000 0 0 $X=11872000 $Y=12624000
X2949 24 2913 buf02 $T=11896000 10072000 0 0 $X=11896000 $Y=10072000
X2950 24 2914 buf02 $T=11937500 12160000 1 180 $X=11904000 $Y=12160000
X2951 24 2915 buf02 $T=11912000 12856000 0 0 $X=11912000 $Y=12856000
X2952 24 2916 buf02 $T=11936000 10072000 0 0 $X=11936000 $Y=10072000
X2953 24 2917 buf02 $T=11977500 12160000 1 180 $X=11944000 $Y=12160000
X2954 24 2918 buf02 $T=11985500 12856000 1 180 $X=11952000 $Y=12856000
X2955 24 2919 buf02 $T=11992000 9840000 0 0 $X=11992000 $Y=9840000
X2956 24 2920 buf02 $T=12025500 12856000 1 180 $X=11992000 $Y=12856000
X2957 24 2921 buf02 $T=12057500 13088000 1 180 $X=12024000 $Y=13088000
X2958 24 2922 buf02 $T=12089500 13552000 1 180 $X=12056000 $Y=13552000
X2959 24 2923 buf02 $T=12097500 13088000 1 180 $X=12064000 $Y=13088000
X2960 24 2924 buf02 $T=12201500 13088000 1 180 $X=12168000 $Y=13088000
X2961 24 2925 buf02 $T=12224000 10072000 0 0 $X=12224000 $Y=10072000
X2962 2926 24 aoi22 $T=280000 4040000 0 0 $X=280000 $Y=4040000
X2963 2927 24 aoi22 $T=377000 3808000 1 180 $X=328000 $Y=3808000
X2964 2928 24 aoi22 $T=376000 2184000 0 0 $X=376000 $Y=2184000
X2965 2929 24 aoi22 $T=449000 6128000 1 180 $X=400000 $Y=6128000
X2966 2930 24 aoi22 $T=489000 7752000 1 180 $X=440000 $Y=7752000
X2967 2931 24 aoi22 $T=513000 5432000 1 180 $X=464000 $Y=5432000
X2968 2932 24 aoi22 $T=528000 4272000 0 0 $X=528000 $Y=4272000
X2969 2933 24 aoi22 $T=536000 3112000 0 0 $X=536000 $Y=3112000
X2970 2934 24 aoi22 $T=585000 7520000 1 180 $X=536000 $Y=7520000
X2971 2935 24 aoi22 $T=609000 3576000 1 180 $X=560000 $Y=3576000
X2972 2936 24 aoi22 $T=641000 5664000 1 180 $X=592000 $Y=5664000
X2973 2937 24 aoi22 $T=641000 7520000 1 180 $X=592000 $Y=7520000
X2974 2938 24 aoi22 $T=665000 3576000 1 180 $X=616000 $Y=3576000
X2975 2939 24 aoi22 $T=673000 11696000 1 180 $X=624000 $Y=11696000
X2976 2940 24 aoi22 $T=648000 7288000 0 0 $X=648000 $Y=7288000
X2977 2941 24 aoi22 $T=697000 11000000 1 180 $X=648000 $Y=11000000
X2978 2942 24 aoi22 $T=697000 11232000 1 180 $X=648000 $Y=11232000
X2979 2943 24 aoi22 $T=729000 6360000 1 180 $X=680000 $Y=6360000
X2980 2944 24 aoi22 $T=753000 96000 1 180 $X=704000 $Y=96000
X2981 2945 24 aoi22 $T=704000 328000 0 0 $X=704000 $Y=328000
X2982 2946 24 aoi22 $T=753000 6128000 1 180 $X=704000 $Y=6128000
X2983 2947 24 aoi22 $T=753000 7520000 1 180 $X=704000 $Y=7520000
X2984 2948 24 aoi22 $T=704000 8216000 0 0 $X=704000 $Y=8216000
X2985 2949 24 aoi22 $T=736000 7752000 0 0 $X=736000 $Y=7752000
X2986 2950 24 aoi22 $T=793000 7056000 1 180 $X=744000 $Y=7056000
X2987 2951 24 aoi22 $T=793000 11928000 1 180 $X=744000 $Y=11928000
X2988 2952 24 aoi22 $T=809000 4736000 1 180 $X=760000 $Y=4736000
X2989 2953 24 aoi22 $T=809000 13088000 1 180 $X=760000 $Y=13088000
X2990 2954 24 aoi22 $T=817000 5432000 1 180 $X=768000 $Y=5432000
X2991 2955 24 aoi22 $T=825000 10072000 1 180 $X=776000 $Y=10072000
X2992 2956 24 aoi22 $T=816000 6128000 0 0 $X=816000 $Y=6128000
X2993 2957 24 aoi22 $T=865000 13088000 1 180 $X=816000 $Y=13088000
X2994 2958 24 aoi22 $T=913000 5200000 1 180 $X=864000 $Y=5200000
X2995 2959 24 aoi22 $T=864000 11464000 0 0 $X=864000 $Y=11464000
X2996 2960 24 aoi22 $T=872000 13320000 0 0 $X=872000 $Y=13320000
X2997 2961 24 aoi22 $T=928000 13320000 0 0 $X=928000 $Y=13320000
X2998 2962 24 aoi22 $T=936000 12856000 0 0 $X=936000 $Y=12856000
X2999 2963 24 aoi22 $T=1033000 560000 1 180 $X=984000 $Y=560000
X3000 2964 24 aoi22 $T=1033000 2648000 1 180 $X=984000 $Y=2648000
X3001 2965 24 aoi22 $T=1041000 5664000 1 180 $X=992000 $Y=5664000
X3002 2966 24 aoi22 $T=1041000 12856000 1 180 $X=992000 $Y=12856000
X3003 2967 24 aoi22 $T=1097000 12856000 1 180 $X=1048000 $Y=12856000
X3004 2968 24 aoi22 $T=1105000 7288000 1 180 $X=1056000 $Y=7288000
X3005 2969 24 aoi22 $T=1113000 9144000 1 180 $X=1064000 $Y=9144000
X3006 2970 24 aoi22 $T=1137000 4504000 1 180 $X=1088000 $Y=4504000
X3007 2971 24 aoi22 $T=1153000 6592000 1 180 $X=1104000 $Y=6592000
X3008 2972 24 aoi22 $T=1153000 7984000 1 180 $X=1104000 $Y=7984000
X3009 2973 24 aoi22 $T=1153000 12856000 1 180 $X=1104000 $Y=12856000
X3010 2974 24 aoi22 $T=1161000 5664000 1 180 $X=1112000 $Y=5664000
X3011 2975 24 aoi22 $T=1161000 7520000 1 180 $X=1112000 $Y=7520000
X3012 2976 24 aoi22 $T=1128000 2184000 0 0 $X=1128000 $Y=2184000
X3013 2977 24 aoi22 $T=1193000 4504000 1 180 $X=1144000 $Y=4504000
X3014 2978 24 aoi22 $T=1168000 7520000 0 0 $X=1168000 $Y=7520000
X3015 2979 24 aoi22 $T=1217000 8448000 1 180 $X=1168000 $Y=8448000
X3016 2980 24 aoi22 $T=1217000 9376000 1 180 $X=1168000 $Y=9376000
X3017 2981 24 aoi22 $T=1225000 9608000 1 180 $X=1176000 $Y=9608000
X3018 2982 24 aoi22 $T=1176000 11464000 0 0 $X=1176000 $Y=11464000
X3019 2983 24 aoi22 $T=1233000 8912000 1 180 $X=1184000 $Y=8912000
X3020 2984 24 aoi22 $T=1241000 1952000 1 180 $X=1192000 $Y=1952000
X3021 2985 24 aoi22 $T=1200000 4504000 0 0 $X=1200000 $Y=4504000
X3022 2986 24 aoi22 $T=1216000 7752000 0 0 $X=1216000 $Y=7752000
X3023 2987 24 aoi22 $T=1216000 12856000 0 0 $X=1216000 $Y=12856000
X3024 2988 24 aoi22 $T=1224000 4968000 0 0 $X=1224000 $Y=4968000
X3025 2989 24 aoi22 $T=1273000 9376000 1 180 $X=1224000 $Y=9376000
X3026 2990 24 aoi22 $T=1232000 792000 0 0 $X=1232000 $Y=792000
X3027 2991 24 aoi22 $T=1232000 6128000 0 0 $X=1232000 $Y=6128000
X3028 2992 24 aoi22 $T=1232000 11928000 0 0 $X=1232000 $Y=11928000
X3029 2993 24 aoi22 $T=1240000 5432000 0 0 $X=1240000 $Y=5432000
X3030 2994 24 aoi22 $T=1289000 8912000 1 180 $X=1240000 $Y=8912000
X3031 2995 24 aoi22 $T=1256000 7984000 0 0 $X=1256000 $Y=7984000
X3032 2996 24 aoi22 $T=1288000 11232000 0 0 $X=1288000 $Y=11232000
X3033 2997 24 aoi22 $T=1296000 8912000 0 0 $X=1296000 $Y=8912000
X3034 2998 24 aoi22 $T=1361000 1256000 1 180 $X=1312000 $Y=1256000
X3035 2999 24 aoi22 $T=1312000 9144000 0 0 $X=1312000 $Y=9144000
X3036 3000 24 aoi22 $T=1384000 13088000 0 0 $X=1384000 $Y=13088000
X3037 3001 24 aoi22 $T=1505000 2880000 1 180 $X=1456000 $Y=2880000
X3038 3002 24 aoi22 $T=1505000 9608000 1 180 $X=1456000 $Y=9608000
X3039 3003 24 aoi22 $T=1513000 12392000 1 180 $X=1464000 $Y=12392000
X3040 3004 24 aoi22 $T=1793000 11000000 1 180 $X=1744000 $Y=11000000
X3041 3005 24 aoi22 $T=1809000 4504000 1 180 $X=1760000 $Y=4504000
X3042 3006 24 aoi22 $T=1825000 4968000 1 180 $X=1776000 $Y=4968000
X3043 3007 24 aoi22 $T=1833000 9376000 1 180 $X=1784000 $Y=9376000
X3044 3008 24 aoi22 $T=1792000 11464000 0 0 $X=1792000 $Y=11464000
X3045 3009 24 aoi22 $T=1873000 12392000 1 180 $X=1824000 $Y=12392000
X3046 3010 24 aoi22 $T=1873000 13320000 1 180 $X=1824000 $Y=13320000
X3047 3011 24 aoi22 $T=1840000 9608000 0 0 $X=1840000 $Y=9608000
X3048 3012 24 aoi22 $T=1897000 4736000 1 180 $X=1848000 $Y=4736000
X3049 3013 24 aoi22 $T=1856000 8216000 0 0 $X=1856000 $Y=8216000
X3050 3014 24 aoi22 $T=1864000 7752000 0 0 $X=1864000 $Y=7752000
X3051 3015 24 aoi22 $T=1913000 10768000 1 180 $X=1864000 $Y=10768000
X3052 3016 24 aoi22 $T=1888000 2416000 0 0 $X=1888000 $Y=2416000
X3053 3017 24 aoi22 $T=1896000 9608000 0 0 $X=1896000 $Y=9608000
X3054 3018 24 aoi22 $T=1953000 6592000 1 180 $X=1904000 $Y=6592000
X3055 3019 24 aoi22 $T=1928000 7288000 0 0 $X=1928000 $Y=7288000
X3056 3020 24 aoi22 $T=1977000 13088000 1 180 $X=1928000 $Y=13088000
X3057 3021 24 aoi22 $T=1976000 12392000 0 0 $X=1976000 $Y=12392000
X3058 3022 24 aoi22 $T=2041000 6128000 1 180 $X=1992000 $Y=6128000
X3059 3023 24 aoi22 $T=2057000 5432000 1 180 $X=2008000 $Y=5432000
X3060 3024 24 aoi22 $T=2016000 7288000 0 0 $X=2016000 $Y=7288000
X3061 3025 24 aoi22 $T=2040000 13088000 0 0 $X=2040000 $Y=13088000
X3062 3026 24 aoi22 $T=2080000 6360000 0 0 $X=2080000 $Y=6360000
X3063 3027 24 aoi22 $T=2161000 4504000 1 180 $X=2112000 $Y=4504000
X3064 3028 24 aoi22 $T=2120000 7984000 0 0 $X=2120000 $Y=7984000
X3065 3029 24 aoi22 $T=2128000 3808000 0 0 $X=2128000 $Y=3808000
X3066 3030 24 aoi22 $T=2136000 1720000 0 0 $X=2136000 $Y=1720000
X3067 3031 24 aoi22 $T=2160000 1488000 0 0 $X=2160000 $Y=1488000
X3068 3032 24 aoi22 $T=2209000 5896000 1 180 $X=2160000 $Y=5896000
X3069 3033 24 aoi22 $T=2216000 5896000 0 0 $X=2216000 $Y=5896000
X3070 3034 24 aoi22 $T=2281000 11000000 1 180 $X=2232000 $Y=11000000
X3071 3035 24 aoi22 $T=2240000 7520000 0 0 $X=2240000 $Y=7520000
X3072 3036 24 aoi22 $T=2240000 8448000 0 0 $X=2240000 $Y=8448000
X3073 3037 24 aoi22 $T=2256000 8912000 0 0 $X=2256000 $Y=8912000
X3074 3038 24 aoi22 $T=2337000 328000 1 180 $X=2288000 $Y=328000
X3075 3039 24 aoi22 $T=2328000 5896000 0 0 $X=2328000 $Y=5896000
X3076 3040 24 aoi22 $T=2352000 13320000 0 0 $X=2352000 $Y=13320000
X3077 2304 24 aoi22 $T=2417000 3576000 1 180 $X=2368000 $Y=3576000
X3078 3041 24 aoi22 $T=2417000 9376000 1 180 $X=2368000 $Y=9376000
X3079 3042 24 aoi22 $T=2433000 12392000 1 180 $X=2384000 $Y=12392000
X3080 3043 24 aoi22 $T=2449000 4736000 1 180 $X=2400000 $Y=4736000
X3081 3044 24 aoi22 $T=2481000 3576000 1 180 $X=2432000 $Y=3576000
X3082 3045 24 aoi22 $T=2432000 11464000 0 0 $X=2432000 $Y=11464000
X3083 3046 24 aoi22 $T=2464000 5664000 0 0 $X=2464000 $Y=5664000
X3084 3047 24 aoi22 $T=2488000 3808000 0 0 $X=2488000 $Y=3808000
X3085 3048 24 aoi22 $T=2545000 9608000 1 180 $X=2496000 $Y=9608000
X3086 3049 24 aoi22 $T=2520000 4736000 0 0 $X=2520000 $Y=4736000
X3087 3050 24 aoi22 $T=2520000 11232000 0 0 $X=2520000 $Y=11232000
X3088 3051 24 aoi22 $T=2528000 10768000 0 0 $X=2528000 $Y=10768000
X3089 3052 24 aoi22 $T=2608000 7984000 0 0 $X=2608000 $Y=7984000
X3090 3053 24 aoi22 $T=2608000 9608000 0 0 $X=2608000 $Y=9608000
X3091 3054 24 aoi22 $T=2657000 12624000 1 180 $X=2608000 $Y=12624000
X3092 3055 24 aoi22 $T=2673000 7288000 1 180 $X=2624000 $Y=7288000
X3093 3056 24 aoi22 $T=2648000 1952000 0 0 $X=2648000 $Y=1952000
X3094 3057 24 aoi22 $T=2664000 9608000 0 0 $X=2664000 $Y=9608000
X3095 3058 24 aoi22 $T=2737000 6128000 1 180 $X=2688000 $Y=6128000
X3096 3059 24 aoi22 $T=2745000 3344000 1 180 $X=2696000 $Y=3344000
X3097 3060 24 aoi22 $T=2696000 6360000 0 0 $X=2696000 $Y=6360000
X3098 3061 24 aoi22 $T=2761000 9376000 1 180 $X=2712000 $Y=9376000
X3099 3062 24 aoi22 $T=2712000 13320000 0 0 $X=2712000 $Y=13320000
X3100 3063 24 aoi22 $T=2736000 7288000 0 0 $X=2736000 $Y=7288000
X3101 3064 24 aoi22 $T=2793000 12856000 1 180 $X=2744000 $Y=12856000
X3102 3065 24 aoi22 $T=2760000 5664000 0 0 $X=2760000 $Y=5664000
X3103 3066 24 aoi22 $T=2776000 96000 0 0 $X=2776000 $Y=96000
X3104 3067 24 aoi22 $T=2833000 9144000 1 180 $X=2784000 $Y=9144000
X3105 3068 24 aoi22 $T=2792000 7288000 0 0 $X=2792000 $Y=7288000
X3106 3069 24 aoi22 $T=2857000 8912000 1 180 $X=2808000 $Y=8912000
X3107 3070 24 aoi22 $T=2865000 5896000 1 180 $X=2816000 $Y=5896000
X3108 3071 24 aoi22 $T=2824000 8448000 0 0 $X=2824000 $Y=8448000
X3109 3072 24 aoi22 $T=2856000 12856000 0 0 $X=2856000 $Y=12856000
X3110 3073 24 aoi22 $T=2872000 13320000 0 0 $X=2872000 $Y=13320000
X3111 3074 24 aoi22 $T=2880000 8448000 0 0 $X=2880000 $Y=8448000
X3112 3075 24 aoi22 $T=2912000 12856000 0 0 $X=2912000 $Y=12856000
X3113 3076 24 aoi22 $T=2928000 4736000 0 0 $X=2928000 $Y=4736000
X3114 3077 24 aoi22 $T=2936000 4504000 0 0 $X=2936000 $Y=4504000
X3115 3078 24 aoi22 $T=2968000 7984000 0 0 $X=2968000 $Y=7984000
X3116 3079 24 aoi22 $T=2984000 1256000 0 0 $X=2984000 $Y=1256000
X3117 3080 24 aoi22 $T=3024000 1024000 0 0 $X=3024000 $Y=1024000
X3118 3081 24 aoi22 $T=3089000 96000 1 180 $X=3040000 $Y=96000
X3119 3082 24 aoi22 $T=3040000 3576000 0 0 $X=3040000 $Y=3576000
X3120 3083 24 aoi22 $T=3072000 1488000 0 0 $X=3072000 $Y=1488000
X3121 3084 24 aoi22 $T=3137000 12392000 1 180 $X=3088000 $Y=12392000
X3122 3085 24 aoi22 $T=3145000 11000000 1 180 $X=3096000 $Y=11000000
X3123 3086 24 aoi22 $T=3112000 3808000 0 0 $X=3112000 $Y=3808000
X3124 3087 24 aoi22 $T=3201000 11000000 1 180 $X=3152000 $Y=11000000
X3125 3088 24 aoi22 $T=3264000 11000000 0 0 $X=3264000 $Y=11000000
X3126 3089 24 aoi22 $T=3345000 10768000 1 180 $X=3296000 $Y=10768000
X3127 3090 24 aoi22 $T=3369000 9144000 1 180 $X=3320000 $Y=9144000
X3128 3091 24 aoi22 $T=3320000 11000000 0 0 $X=3320000 $Y=11000000
X3129 3092 24 aoi22 $T=3377000 11464000 1 180 $X=3328000 $Y=11464000
X3130 3093 24 aoi22 $T=3377000 12160000 1 180 $X=3328000 $Y=12160000
X3131 3094 24 aoi22 $T=3376000 12856000 0 0 $X=3376000 $Y=12856000
X3132 3095 24 aoi22 $T=3441000 6592000 1 180 $X=3392000 $Y=6592000
X3133 3096 24 aoi22 $T=3457000 11464000 1 180 $X=3408000 $Y=11464000
X3134 3097 24 aoi22 $T=3481000 9144000 1 180 $X=3432000 $Y=9144000
X3135 3098 24 aoi22 $T=3440000 12392000 0 0 $X=3440000 $Y=12392000
X3136 3099 24 aoi22 $T=3497000 10768000 1 180 $X=3448000 $Y=10768000
X3137 3100 24 aoi22 $T=3545000 8912000 1 180 $X=3496000 $Y=8912000
X3138 3101 24 aoi22 $T=3553000 8680000 1 180 $X=3504000 $Y=8680000
X3139 3102 24 aoi22 $T=3553000 10768000 1 180 $X=3504000 $Y=10768000
X3140 3103 24 aoi22 $T=3520000 11464000 0 0 $X=3520000 $Y=11464000
X3141 3104 24 aoi22 $T=3568000 9840000 0 0 $X=3568000 $Y=9840000
X3142 3105 24 aoi22 $T=3576000 9608000 0 0 $X=3576000 $Y=9608000
X3143 3106 24 aoi22 $T=3665000 5432000 1 180 $X=3616000 $Y=5432000
X3144 3107 24 aoi22 $T=3616000 10768000 0 0 $X=3616000 $Y=10768000
X3145 3108 24 aoi22 $T=3673000 2648000 1 180 $X=3624000 $Y=2648000
X3146 3109 24 aoi22 $T=3624000 11000000 0 0 $X=3624000 $Y=11000000
X3147 3110 24 aoi22 $T=3648000 328000 0 0 $X=3648000 $Y=328000
X3148 3111 24 aoi22 $T=3697000 4040000 1 180 $X=3648000 $Y=4040000
X3149 3112 24 aoi22 $T=3648000 7752000 0 0 $X=3648000 $Y=7752000
X3150 3113 24 aoi22 $T=3705000 7520000 1 180 $X=3656000 $Y=7520000
X3151 3114 24 aoi22 $T=3721000 2880000 1 180 $X=3672000 $Y=2880000
X3152 3115 24 aoi22 $T=3721000 5200000 1 180 $X=3672000 $Y=5200000
X3153 3116 24 aoi22 $T=3672000 11232000 0 0 $X=3672000 $Y=11232000
X3154 3117 24 aoi22 $T=3729000 6360000 1 180 $X=3680000 $Y=6360000
X3155 3118 24 aoi22 $T=3737000 11928000 1 180 $X=3688000 $Y=11928000
X3156 3119 24 aoi22 $T=3745000 2416000 1 180 $X=3696000 $Y=2416000
X3157 3120 24 aoi22 $T=3753000 7752000 1 180 $X=3704000 $Y=7752000
X3158 3121 24 aoi22 $T=3777000 4968000 1 180 $X=3728000 $Y=4968000
X3159 3122 24 aoi22 $T=3728000 5432000 0 0 $X=3728000 $Y=5432000
X3160 3123 24 aoi22 $T=3777000 7288000 1 180 $X=3728000 $Y=7288000
X3161 3124 24 aoi22 $T=3736000 96000 0 0 $X=3736000 $Y=96000
X3162 3125 24 aoi22 $T=3744000 9376000 0 0 $X=3744000 $Y=9376000
X3163 3126 24 aoi22 $T=3760000 6128000 0 0 $X=3760000 $Y=6128000
X3164 3127 24 aoi22 $T=3817000 792000 1 180 $X=3768000 $Y=792000
X3165 3128 24 aoi22 $T=3784000 5432000 0 0 $X=3784000 $Y=5432000
X3166 3129 24 aoi22 $T=3800000 5896000 0 0 $X=3800000 $Y=5896000
X3167 3130 24 aoi22 $T=3873000 792000 1 180 $X=3824000 $Y=792000
X3168 3131 24 aoi22 $T=3832000 9144000 0 0 $X=3832000 $Y=9144000
X3169 3132 24 aoi22 $T=3848000 4504000 0 0 $X=3848000 $Y=4504000
X3170 3133 24 aoi22 $T=3856000 4736000 0 0 $X=3856000 $Y=4736000
X3171 3134 24 aoi22 $T=3929000 792000 1 180 $X=3880000 $Y=792000
X3172 3135 24 aoi22 $T=3888000 9144000 0 0 $X=3888000 $Y=9144000
X3173 3136 24 aoi22 $T=3920000 7752000 0 0 $X=3920000 $Y=7752000
X3174 3137 24 aoi22 $T=3944000 12392000 0 0 $X=3944000 $Y=12392000
X3175 3138 24 aoi22 $T=3976000 7752000 0 0 $X=3976000 $Y=7752000
X3176 3139 24 aoi22 $T=3984000 4272000 0 0 $X=3984000 $Y=4272000
X3177 3140 24 aoi22 $T=4041000 12856000 1 180 $X=3992000 $Y=12856000
X3178 3141 24 aoi22 $T=4065000 3576000 1 180 $X=4016000 $Y=3576000
X3179 3142 24 aoi22 $T=4032000 2880000 0 0 $X=4032000 $Y=2880000
X3180 3143 24 aoi22 $T=4056000 12392000 0 0 $X=4056000 $Y=12392000
X3181 3144 24 aoi22 $T=4080000 1952000 0 0 $X=4080000 $Y=1952000
X3182 3145 24 aoi22 $T=4088000 2880000 0 0 $X=4088000 $Y=2880000
X3183 3146 24 aoi22 $T=4088000 12856000 0 0 $X=4088000 $Y=12856000
X3184 3147 24 aoi22 $T=4104000 7056000 0 0 $X=4104000 $Y=7056000
X3185 3148 24 aoi22 $T=4104000 11696000 0 0 $X=4104000 $Y=11696000
X3186 3149 24 aoi22 $T=4112000 8216000 0 0 $X=4112000 $Y=8216000
X3187 3150 24 aoi22 $T=4169000 1256000 1 180 $X=4120000 $Y=1256000
X3188 3151 24 aoi22 $T=4217000 11000000 1 180 $X=4168000 $Y=11000000
X3189 3152 24 aoi22 $T=4176000 96000 0 0 $X=4176000 $Y=96000
X3190 3153 24 aoi22 $T=4240000 1256000 0 0 $X=4240000 $Y=1256000
X3191 3154 24 aoi22 $T=4297000 9840000 1 180 $X=4248000 $Y=9840000
X3192 3155 24 aoi22 $T=4305000 3344000 1 180 $X=4256000 $Y=3344000
X3193 3156 24 aoi22 $T=4256000 7984000 0 0 $X=4256000 $Y=7984000
X3194 3157 24 aoi22 $T=4313000 9376000 1 180 $X=4264000 $Y=9376000
X3195 3158 24 aoi22 $T=4321000 8912000 1 180 $X=4272000 $Y=8912000
X3196 3159 24 aoi22 $T=4280000 1024000 0 0 $X=4280000 $Y=1024000
X3197 3160 24 aoi22 $T=4280000 11000000 0 0 $X=4280000 $Y=11000000
X3198 3161 24 aoi22 $T=4296000 792000 0 0 $X=4296000 $Y=792000
X3199 3162 24 aoi22 $T=4336000 1024000 0 0 $X=4336000 $Y=1024000
X3200 3163 24 aoi22 $T=4385000 2416000 1 180 $X=4336000 $Y=2416000
X3201 3164 24 aoi22 $T=4336000 9840000 0 0 $X=4336000 $Y=9840000
X3202 3165 24 aoi22 $T=4344000 4968000 0 0 $X=4344000 $Y=4968000
X3203 3166 24 aoi22 $T=4401000 5664000 1 180 $X=4352000 $Y=5664000
X3204 3167 24 aoi22 $T=4376000 3344000 0 0 $X=4376000 $Y=3344000
X3205 3168 24 aoi22 $T=4376000 3576000 0 0 $X=4376000 $Y=3576000
X3206 3169 24 aoi22 $T=4376000 9144000 0 0 $X=4376000 $Y=9144000
X3207 3170 24 aoi22 $T=4384000 6128000 0 0 $X=4384000 $Y=6128000
X3208 3171 24 aoi22 $T=4384000 9608000 0 0 $X=4384000 $Y=9608000
X3209 3172 24 aoi22 $T=4392000 3808000 0 0 $X=4392000 $Y=3808000
X3210 3173 24 aoi22 $T=4449000 5432000 1 180 $X=4400000 $Y=5432000
X3211 3174 24 aoi22 $T=4408000 6360000 0 0 $X=4408000 $Y=6360000
X3212 3175 24 aoi22 $T=4416000 10768000 0 0 $X=4416000 $Y=10768000
X3213 3176 24 aoi22 $T=4416000 13088000 0 0 $X=4416000 $Y=13088000
X3214 3177 24 aoi22 $T=4489000 4736000 1 180 $X=4440000 $Y=4736000
X3215 3178 24 aoi22 $T=4440000 9608000 0 0 $X=4440000 $Y=9608000
X3216 3179 24 aoi22 $T=4456000 1024000 0 0 $X=4456000 $Y=1024000
X3217 3180 24 aoi22 $T=4464000 4504000 0 0 $X=4464000 $Y=4504000
X3218 3181 24 aoi22 $T=4480000 12856000 0 0 $X=4480000 $Y=12856000
X3219 3182 24 aoi22 $T=4504000 9144000 0 0 $X=4504000 $Y=9144000
X3220 3183 24 aoi22 $T=4577000 2416000 1 180 $X=4528000 $Y=2416000
X3221 3184 24 aoi22 $T=4608000 2184000 0 0 $X=4608000 $Y=2184000
X3222 3185 24 aoi22 $T=4640000 11464000 0 0 $X=4640000 $Y=11464000
X3223 3186 24 aoi22 $T=4713000 7520000 1 180 $X=4664000 $Y=7520000
X3224 3187 24 aoi22 $T=4696000 11000000 0 0 $X=4696000 $Y=11000000
X3225 3188 24 aoi22 $T=4753000 5432000 1 180 $X=4704000 $Y=5432000
X3226 3189 24 aoi22 $T=4801000 12392000 1 180 $X=4752000 $Y=12392000
X3227 3190 24 aoi22 $T=4760000 5432000 0 0 $X=4760000 $Y=5432000
X3228 3191 24 aoi22 $T=4784000 5896000 0 0 $X=4784000 $Y=5896000
X3229 3192 24 aoi22 $T=4832000 4736000 0 0 $X=4832000 $Y=4736000
X3230 3193 24 aoi22 $T=4840000 5896000 0 0 $X=4840000 $Y=5896000
X3231 3194 24 aoi22 $T=4864000 12392000 0 0 $X=4864000 $Y=12392000
X3232 3195 24 aoi22 $T=4888000 4736000 0 0 $X=4888000 $Y=4736000
X3233 3196 24 aoi22 $T=4896000 5896000 0 0 $X=4896000 $Y=5896000
X3234 3197 24 aoi22 $T=4945000 8448000 1 180 $X=4896000 $Y=8448000
X3235 3198 24 aoi22 $T=4936000 5432000 0 0 $X=4936000 $Y=5432000
X3236 3199 24 aoi22 $T=4952000 5664000 0 0 $X=4952000 $Y=5664000
X3237 3200 24 aoi22 $T=4952000 5896000 0 0 $X=4952000 $Y=5896000
X3238 3201 24 aoi22 $T=4960000 12624000 0 0 $X=4960000 $Y=12624000
X3239 3202 24 aoi22 $T=5025000 9376000 1 180 $X=4976000 $Y=9376000
X3240 3203 24 aoi22 $T=5008000 6128000 0 0 $X=5008000 $Y=6128000
X3241 3204 24 aoi22 $T=5089000 1024000 1 180 $X=5040000 $Y=1024000
X3242 3205 24 aoi22 $T=5048000 792000 0 0 $X=5048000 $Y=792000
X3243 3206 24 aoi22 $T=5056000 5432000 0 0 $X=5056000 $Y=5432000
X3244 3207 24 aoi22 $T=5056000 11000000 0 0 $X=5056000 $Y=11000000
X3245 3208 24 aoi22 $T=5064000 6128000 0 0 $X=5064000 $Y=6128000
X3246 3209 24 aoi22 $T=5121000 7752000 1 180 $X=5072000 $Y=7752000
X3247 3210 24 aoi22 $T=5072000 8680000 0 0 $X=5072000 $Y=8680000
X3248 3211 24 aoi22 $T=5088000 328000 0 0 $X=5088000 $Y=328000
X3249 3212 24 aoi22 $T=5096000 1024000 0 0 $X=5096000 $Y=1024000
X3250 3213 24 aoi22 $T=5153000 2416000 1 180 $X=5104000 $Y=2416000
X3251 3214 24 aoi22 $T=5161000 8216000 1 180 $X=5112000 $Y=8216000
X3252 3215 24 aoi22 $T=5169000 560000 1 180 $X=5120000 $Y=560000
X3253 3216 24 aoi22 $T=5128000 7752000 0 0 $X=5128000 $Y=7752000
X3254 3217 24 aoi22 $T=5193000 328000 1 180 $X=5144000 $Y=328000
X3255 3218 24 aoi22 $T=5152000 6360000 0 0 $X=5152000 $Y=6360000
X3256 3219 24 aoi22 $T=5160000 792000 0 0 $X=5160000 $Y=792000
X3257 3220 24 aoi22 $T=5160000 2416000 0 0 $X=5160000 $Y=2416000
X3258 3221 24 aoi22 $T=5209000 12856000 1 180 $X=5160000 $Y=12856000
X3259 3222 24 aoi22 $T=5184000 11696000 0 0 $X=5184000 $Y=11696000
X3260 3223 24 aoi22 $T=5241000 2880000 1 180 $X=5192000 $Y=2880000
X3261 3224 24 aoi22 $T=5192000 11464000 0 0 $X=5192000 $Y=11464000
X3262 3225 24 aoi22 $T=5208000 8912000 0 0 $X=5208000 $Y=8912000
X3263 3226 24 aoi22 $T=5265000 2416000 1 180 $X=5216000 $Y=2416000
X3264 3227 24 aoi22 $T=5281000 560000 1 180 $X=5232000 $Y=560000
X3265 3228 24 aoi22 $T=5240000 11928000 0 0 $X=5240000 $Y=11928000
X3266 3229 24 aoi22 $T=5297000 2880000 1 180 $X=5248000 $Y=2880000
X3267 3230 24 aoi22 $T=5264000 8912000 0 0 $X=5264000 $Y=8912000
X3268 3231 24 aoi22 $T=5272000 12856000 0 0 $X=5272000 $Y=12856000
X3269 3232 24 aoi22 $T=5280000 9840000 0 0 $X=5280000 $Y=9840000
X3270 3233 24 aoi22 $T=5337000 3112000 1 180 $X=5288000 $Y=3112000
X3271 3234 24 aoi22 $T=5296000 10768000 0 0 $X=5296000 $Y=10768000
X3272 3235 24 aoi22 $T=5312000 2648000 0 0 $X=5312000 $Y=2648000
X3273 3236 24 aoi22 $T=5320000 8912000 0 0 $X=5320000 $Y=8912000
X3274 3237 24 aoi22 $T=5336000 2416000 0 0 $X=5336000 $Y=2416000
X3275 3238 24 aoi22 $T=5336000 11928000 0 0 $X=5336000 $Y=11928000
X3276 3239 24 aoi22 $T=5401000 3344000 1 180 $X=5352000 $Y=3344000
X3277 3240 24 aoi22 $T=5417000 5664000 1 180 $X=5368000 $Y=5664000
X3278 3241 24 aoi22 $T=5384000 560000 0 0 $X=5384000 $Y=560000
X3279 3242 24 aoi22 $T=5392000 4040000 0 0 $X=5392000 $Y=4040000
X3280 3243 24 aoi22 $T=5457000 3344000 1 180 $X=5408000 $Y=3344000
X3281 3244 24 aoi22 $T=5473000 5664000 1 180 $X=5424000 $Y=5664000
X3282 3245 24 aoi22 $T=5432000 9608000 0 0 $X=5432000 $Y=9608000
X3283 3246 24 aoi22 $T=5440000 560000 0 0 $X=5440000 $Y=560000
X3284 3247 24 aoi22 $T=5456000 6360000 0 0 $X=5456000 $Y=6360000
X3285 3248 24 aoi22 $T=5456000 13320000 0 0 $X=5456000 $Y=13320000
X3286 3249 24 aoi22 $T=5480000 6592000 0 0 $X=5480000 $Y=6592000
X3287 3250 24 aoi22 $T=5537000 7752000 1 180 $X=5488000 $Y=7752000
X3288 3251 24 aoi22 $T=5512000 6824000 0 0 $X=5512000 $Y=6824000
X3289 3252 24 aoi22 $T=5569000 7056000 1 180 $X=5520000 $Y=7056000
X3290 3253 24 aoi22 $T=5528000 3808000 0 0 $X=5528000 $Y=3808000
X3291 3254 24 aoi22 $T=5536000 5664000 0 0 $X=5536000 $Y=5664000
X3292 3255 24 aoi22 $T=5544000 7752000 0 0 $X=5544000 $Y=7752000
X3293 3256 24 aoi22 $T=5576000 4736000 0 0 $X=5576000 $Y=4736000
X3294 3257 24 aoi22 $T=5576000 7056000 0 0 $X=5576000 $Y=7056000
X3295 3258 24 aoi22 $T=5633000 2880000 1 180 $X=5584000 $Y=2880000
X3296 3259 24 aoi22 $T=5584000 3808000 0 0 $X=5584000 $Y=3808000
X3297 3260 24 aoi22 $T=5592000 6592000 0 0 $X=5592000 $Y=6592000
X3298 3261 24 aoi22 $T=5616000 2184000 0 0 $X=5616000 $Y=2184000
X3299 3262 24 aoi22 $T=5632000 7752000 0 0 $X=5632000 $Y=7752000
X3300 3263 24 aoi22 $T=5640000 12856000 0 0 $X=5640000 $Y=12856000
X3301 3264 24 aoi22 $T=5697000 12392000 1 180 $X=5648000 $Y=12392000
X3302 3265 24 aoi22 $T=5672000 2184000 0 0 $X=5672000 $Y=2184000
X3303 3266 24 aoi22 $T=5696000 10768000 0 0 $X=5696000 $Y=10768000
X3304 3267 24 aoi22 $T=5801000 328000 1 180 $X=5752000 $Y=328000
X3305 3268 24 aoi22 $T=5801000 9840000 1 180 $X=5752000 $Y=9840000
X3306 3269 24 aoi22 $T=5800000 12624000 0 0 $X=5800000 $Y=12624000
X3307 3270 24 aoi22 $T=5808000 328000 0 0 $X=5808000 $Y=328000
X3308 3271 24 aoi22 $T=5840000 5664000 0 0 $X=5840000 $Y=5664000
X3309 3272 24 aoi22 $T=5913000 2648000 1 180 $X=5864000 $Y=2648000
X3310 3273 24 aoi22 $T=5921000 11696000 1 180 $X=5872000 $Y=11696000
X3311 3274 24 aoi22 $T=5929000 2416000 1 180 $X=5880000 $Y=2416000
X3312 3275 24 aoi22 $T=5888000 7288000 0 0 $X=5888000 $Y=7288000
X3313 3276 24 aoi22 $T=5904000 8912000 0 0 $X=5904000 $Y=8912000
X3314 3277 24 aoi22 $T=5912000 4736000 0 0 $X=5912000 $Y=4736000
X3315 3278 24 aoi22 $T=5969000 1024000 1 180 $X=5920000 $Y=1024000
X3316 3279 24 aoi22 $T=6009000 3344000 1 180 $X=5960000 $Y=3344000
X3317 3280 24 aoi22 $T=6009000 4040000 1 180 $X=5960000 $Y=4040000
X3318 3281 24 aoi22 $T=5968000 7984000 0 0 $X=5968000 $Y=7984000
X3319 3282 24 aoi22 $T=6017000 8680000 1 180 $X=5968000 $Y=8680000
X3320 3283 24 aoi22 $T=6025000 1024000 1 180 $X=5976000 $Y=1024000
X3321 3284 24 aoi22 $T=5976000 2880000 0 0 $X=5976000 $Y=2880000
X3322 3285 24 aoi22 $T=5976000 13320000 0 0 $X=5976000 $Y=13320000
X3323 3286 24 aoi22 $T=6033000 3808000 1 180 $X=5984000 $Y=3808000
X3324 3287 24 aoi22 $T=5984000 11696000 0 0 $X=5984000 $Y=11696000
X3325 3288 24 aoi22 $T=5992000 2416000 0 0 $X=5992000 $Y=2416000
X3326 3289 24 aoi22 $T=5992000 10768000 0 0 $X=5992000 $Y=10768000
X3327 3290 24 aoi22 $T=5992000 11928000 0 0 $X=5992000 $Y=11928000
X3328 3291 24 aoi22 $T=5992000 12856000 0 0 $X=5992000 $Y=12856000
X3329 3292 24 aoi22 $T=6000000 11000000 0 0 $X=6000000 $Y=11000000
X3330 3293 24 aoi22 $T=6008000 7288000 0 0 $X=6008000 $Y=7288000
X3331 3294 24 aoi22 $T=6024000 792000 0 0 $X=6024000 $Y=792000
X3332 3295 24 aoi22 $T=6024000 12392000 0 0 $X=6024000 $Y=12392000
X3333 3296 24 aoi22 $T=6089000 3808000 1 180 $X=6040000 $Y=3808000
X3334 3297 24 aoi22 $T=6040000 12624000 0 0 $X=6040000 $Y=12624000
X3335 3298 24 aoi22 $T=6056000 7752000 0 0 $X=6056000 $Y=7752000
X3336 3299 24 aoi22 $T=6088000 9608000 0 0 $X=6088000 $Y=9608000
X3337 3300 24 aoi22 $T=6112000 2416000 0 0 $X=6112000 $Y=2416000
X3338 3301 24 aoi22 $T=6152000 3808000 0 0 $X=6152000 $Y=3808000
X3339 3302 24 aoi22 $T=6320000 3344000 0 0 $X=6320000 $Y=3344000
X3340 3303 24 aoi22 $T=6441000 5432000 1 180 $X=6392000 $Y=5432000
X3341 3304 24 aoi22 $T=6441000 6128000 1 180 $X=6392000 $Y=6128000
X3342 3305 24 aoi22 $T=6545000 328000 1 180 $X=6496000 $Y=328000
X3343 3306 24 aoi22 $T=6641000 2880000 1 180 $X=6592000 $Y=2880000
X3344 3307 24 aoi22 $T=6641000 6824000 1 180 $X=6592000 $Y=6824000
X3345 3308 24 aoi22 $T=6616000 4504000 0 0 $X=6616000 $Y=4504000
X3346 3309 24 aoi22 $T=6681000 6592000 1 180 $X=6632000 $Y=6592000
X3347 3310 24 aoi22 $T=6729000 1024000 1 180 $X=6680000 $Y=1024000
X3348 3311 24 aoi22 $T=6737000 2416000 1 180 $X=6688000 $Y=2416000
X3349 3312 24 aoi22 $T=6688000 3576000 0 0 $X=6688000 $Y=3576000
X3350 3313 24 aoi22 $T=6712000 3112000 0 0 $X=6712000 $Y=3112000
X3351 3314 24 aoi22 $T=6769000 1952000 1 180 $X=6720000 $Y=1952000
X3352 3315 24 aoi22 $T=6720000 6128000 0 0 $X=6720000 $Y=6128000
X3353 3316 24 aoi22 $T=6769000 10536000 1 180 $X=6720000 $Y=10536000
X3354 3317 24 aoi22 $T=6785000 1024000 1 180 $X=6736000 $Y=1024000
X3355 3318 24 aoi22 $T=6744000 3576000 0 0 $X=6744000 $Y=3576000
X3356 3319 24 aoi22 $T=6801000 9376000 1 180 $X=6752000 $Y=9376000
X3357 3320 24 aoi22 $T=6768000 2880000 0 0 $X=6768000 $Y=2880000
X3358 3321 24 aoi22 $T=6776000 6128000 0 0 $X=6776000 $Y=6128000
X3359 3322 24 aoi22 $T=6825000 10536000 1 180 $X=6776000 $Y=10536000
X3360 3323 24 aoi22 $T=6833000 12392000 1 180 $X=6784000 $Y=12392000
X3361 3324 24 aoi22 $T=6849000 13088000 1 180 $X=6800000 $Y=13088000
X3362 3325 24 aoi22 $T=6848000 11464000 0 0 $X=6848000 $Y=11464000
X3363 3326 24 aoi22 $T=6905000 13088000 1 180 $X=6856000 $Y=13088000
X3364 3327 24 aoi22 $T=6872000 2184000 0 0 $X=6872000 $Y=2184000
X3365 3328 24 aoi22 $T=6929000 11232000 1 180 $X=6880000 $Y=11232000
X3366 3329 24 aoi22 $T=6888000 6128000 0 0 $X=6888000 $Y=6128000
X3367 3330 24 aoi22 $T=6888000 8912000 0 0 $X=6888000 $Y=8912000
X3368 3331 24 aoi22 $T=6888000 11696000 0 0 $X=6888000 $Y=11696000
X3369 3332 24 aoi22 $T=6985000 9840000 1 180 $X=6936000 $Y=9840000
X3370 3333 24 aoi22 $T=6944000 6128000 0 0 $X=6944000 $Y=6128000
X3371 3334 24 aoi22 $T=6944000 11696000 0 0 $X=6944000 $Y=11696000
X3372 3335 24 aoi22 $T=6960000 11000000 0 0 $X=6960000 $Y=11000000
X3373 3336 24 aoi22 $T=6968000 792000 0 0 $X=6968000 $Y=792000
X3374 3337 24 aoi22 $T=6976000 560000 0 0 $X=6976000 $Y=560000
X3375 3338 24 aoi22 $T=7025000 9144000 1 180 $X=6976000 $Y=9144000
X3376 3339 24 aoi22 $T=6984000 4272000 0 0 $X=6984000 $Y=4272000
X3377 3340 24 aoi22 $T=6992000 8912000 0 0 $X=6992000 $Y=8912000
X3378 3341 24 aoi22 $T=7000000 11464000 0 0 $X=7000000 $Y=11464000
X3379 3342 24 aoi22 $T=7024000 2648000 0 0 $X=7024000 $Y=2648000
X3380 3343 24 aoi22 $T=7048000 9840000 0 0 $X=7048000 $Y=9840000
X3381 3344 24 aoi22 $T=7105000 13552000 1 180 $X=7056000 $Y=13552000
X3382 3345 24 aoi22 $T=7080000 10536000 0 0 $X=7080000 $Y=10536000
X3383 3346 24 aoi22 $T=7153000 3576000 1 180 $X=7104000 $Y=3576000
X3384 3347 24 aoi22 $T=7177000 7520000 1 180 $X=7128000 $Y=7520000
X3385 3348 24 aoi22 $T=7136000 9376000 0 0 $X=7136000 $Y=9376000
X3386 3349 24 aoi22 $T=7233000 7520000 1 180 $X=7184000 $Y=7520000
X3387 3350 24 aoi22 $T=7184000 12856000 0 0 $X=7184000 $Y=12856000
X3388 3351 24 aoi22 $T=7224000 4736000 0 0 $X=7224000 $Y=4736000
X3389 3352 24 aoi22 $T=7289000 7520000 1 180 $X=7240000 $Y=7520000
X3390 3353 24 aoi22 $T=7272000 1256000 0 0 $X=7272000 $Y=1256000
X3391 3354 24 aoi22 $T=7272000 3808000 0 0 $X=7272000 $Y=3808000
X3392 3355 24 aoi22 $T=7280000 4504000 0 0 $X=7280000 $Y=4504000
X3393 3356 24 aoi22 $T=7345000 7984000 1 180 $X=7296000 $Y=7984000
X3394 3357 24 aoi22 $T=7328000 1952000 0 0 $X=7328000 $Y=1952000
X3395 3358 24 aoi22 $T=7328000 3344000 0 0 $X=7328000 $Y=3344000
X3396 3359 24 aoi22 $T=7328000 3808000 0 0 $X=7328000 $Y=3808000
X3397 3360 24 aoi22 $T=7352000 7520000 0 0 $X=7352000 $Y=7520000
X3398 3361 24 aoi22 $T=7400000 12624000 0 0 $X=7400000 $Y=12624000
X3399 3362 24 aoi22 $T=7408000 4040000 0 0 $X=7408000 $Y=4040000
X3400 3363 24 aoi22 $T=7408000 7288000 0 0 $X=7408000 $Y=7288000
X3401 3364 24 aoi22 $T=7408000 12392000 0 0 $X=7408000 $Y=12392000
X3402 3365 24 aoi22 $T=7424000 2184000 0 0 $X=7424000 $Y=2184000
X3403 3366 24 aoi22 $T=7440000 4504000 0 0 $X=7440000 $Y=4504000
X3404 3367 24 aoi22 $T=7505000 5664000 1 180 $X=7456000 $Y=5664000
X3405 3368 24 aoi22 $T=7529000 8216000 1 180 $X=7480000 $Y=8216000
X3406 3369 24 aoi22 $T=7480000 8912000 0 0 $X=7480000 $Y=8912000
X3407 3370 24 aoi22 $T=7561000 5664000 1 180 $X=7512000 $Y=5664000
X3408 3371 24 aoi22 $T=7512000 13088000 0 0 $X=7512000 $Y=13088000
X3409 3372 24 aoi22 $T=7528000 1024000 0 0 $X=7528000 $Y=1024000
X3410 3373 24 aoi22 $T=7585000 8912000 1 180 $X=7536000 $Y=8912000
X3411 3374 24 aoi22 $T=7617000 5664000 1 180 $X=7568000 $Y=5664000
X3412 3375 24 aoi22 $T=7568000 13088000 0 0 $X=7568000 $Y=13088000
X3413 3376 24 aoi22 $T=7576000 2648000 0 0 $X=7576000 $Y=2648000
X3414 3377 24 aoi22 $T=7584000 1024000 0 0 $X=7584000 $Y=1024000
X3415 3378 24 aoi22 $T=7592000 13320000 0 0 $X=7592000 $Y=13320000
X3416 3379 24 aoi22 $T=7616000 2880000 0 0 $X=7616000 $Y=2880000
X3417 3380 24 aoi22 $T=7648000 7984000 0 0 $X=7648000 $Y=7984000
X3418 3381 24 aoi22 $T=7648000 8912000 0 0 $X=7648000 $Y=8912000
X3419 3382 24 aoi22 $T=7697000 11696000 1 180 $X=7648000 $Y=11696000
X3420 3383 24 aoi22 $T=7656000 7520000 0 0 $X=7656000 $Y=7520000
X3421 3384 24 aoi22 $T=7680000 5664000 0 0 $X=7680000 $Y=5664000
X3422 3385 24 aoi22 $T=7745000 10304000 1 180 $X=7696000 $Y=10304000
X3423 3386 24 aoi22 $T=7801000 10304000 1 180 $X=7752000 $Y=10304000
X3424 3387 24 aoi22 $T=7792000 5664000 0 0 $X=7792000 $Y=5664000
X3425 3388 24 aoi22 $T=7824000 5432000 0 0 $X=7824000 $Y=5432000
X3426 3389 24 aoi22 $T=7921000 560000 1 180 $X=7872000 $Y=560000
X3427 3390 24 aoi22 $T=7969000 7984000 1 180 $X=7920000 $Y=7984000
X3428 3391 24 aoi22 $T=7993000 2416000 1 180 $X=7944000 $Y=2416000
X3429 3392 24 aoi22 $T=8009000 7520000 1 180 $X=7960000 $Y=7520000
X3430 3393 24 aoi22 $T=8025000 7984000 1 180 $X=7976000 $Y=7984000
X3431 3394 24 aoi22 $T=8016000 12392000 0 0 $X=8016000 $Y=12392000
X3432 3395 24 aoi22 $T=8024000 7288000 0 0 $X=8024000 $Y=7288000
X3433 3396 24 aoi22 $T=8113000 7752000 1 180 $X=8064000 $Y=7752000
X3434 3397 24 aoi22 $T=8072000 7520000 0 0 $X=8072000 $Y=7520000
X3435 3398 24 aoi22 $T=8072000 12392000 0 0 $X=8072000 $Y=12392000
X3436 3399 24 aoi22 $T=8137000 11696000 1 180 $X=8088000 $Y=11696000
X3437 3400 24 aoi22 $T=8145000 1720000 1 180 $X=8096000 $Y=1720000
X3438 3401 24 aoi22 $T=8096000 5664000 0 0 $X=8096000 $Y=5664000
X3439 3402 24 aoi22 $T=8153000 792000 1 180 $X=8104000 $Y=792000
X3440 3403 24 aoi22 $T=8112000 1952000 0 0 $X=8112000 $Y=1952000
X3441 3404 24 aoi22 $T=8177000 10304000 1 180 $X=8128000 $Y=10304000
X3442 3405 24 aoi22 $T=8136000 2880000 0 0 $X=8136000 $Y=2880000
X3443 3406 24 aoi22 $T=8209000 792000 1 180 $X=8160000 $Y=792000
X3444 3407 24 aoi22 $T=8209000 3808000 1 180 $X=8160000 $Y=3808000
X3445 3408 24 aoi22 $T=8209000 9840000 1 180 $X=8160000 $Y=9840000
X3446 3409 24 aoi22 $T=8168000 1952000 0 0 $X=8168000 $Y=1952000
X3447 3410 24 aoi22 $T=8184000 12392000 0 0 $X=8184000 $Y=12392000
X3448 3411 24 aoi22 $T=8192000 2880000 0 0 $X=8192000 $Y=2880000
X3449 3412 24 aoi22 $T=8200000 11696000 0 0 $X=8200000 $Y=11696000
X3450 3413 24 aoi22 $T=8208000 5664000 0 0 $X=8208000 $Y=5664000
X3451 3414 24 aoi22 $T=8265000 9840000 1 180 $X=8216000 $Y=9840000
X3452 3415 24 aoi22 $T=8264000 5664000 0 0 $X=8264000 $Y=5664000
X3453 3416 24 aoi22 $T=8280000 2416000 0 0 $X=8280000 $Y=2416000
X3454 3417 24 aoi22 $T=8296000 12392000 0 0 $X=8296000 $Y=12392000
X3455 3418 24 aoi22 $T=8304000 792000 0 0 $X=8304000 $Y=792000
X3456 3419 24 aoi22 $T=8304000 3808000 0 0 $X=8304000 $Y=3808000
X3457 3420 24 aoi22 $T=8353000 13320000 1 180 $X=8304000 $Y=13320000
X3458 3421 24 aoi22 $T=8369000 6128000 1 180 $X=8320000 $Y=6128000
X3459 3422 24 aoi22 $T=8320000 10072000 0 0 $X=8320000 $Y=10072000
X3460 3423 24 aoi22 $T=8328000 1952000 0 0 $X=8328000 $Y=1952000
X3461 3424 24 aoi22 $T=8377000 8912000 1 180 $X=8328000 $Y=8912000
X3462 3425 24 aoi22 $T=8336000 2416000 0 0 $X=8336000 $Y=2416000
X3463 3426 24 aoi22 $T=8352000 2880000 0 0 $X=8352000 $Y=2880000
X3464 3427 24 aoi22 $T=8352000 12392000 0 0 $X=8352000 $Y=12392000
X3465 3428 24 aoi22 $T=8360000 13320000 0 0 $X=8360000 $Y=13320000
X3466 3429 24 aoi22 $T=8417000 6360000 1 180 $X=8368000 $Y=6360000
X3467 3430 24 aoi22 $T=8441000 328000 1 180 $X=8392000 $Y=328000
X3468 3431 24 aoi22 $T=8408000 2880000 0 0 $X=8408000 $Y=2880000
X3469 3432 24 aoi22 $T=8408000 12392000 0 0 $X=8408000 $Y=12392000
X3470 3433 24 aoi22 $T=8424000 3808000 0 0 $X=8424000 $Y=3808000
X3471 3434 24 aoi22 $T=8505000 4504000 1 180 $X=8456000 $Y=4504000
X3472 3435 24 aoi22 $T=8456000 9376000 0 0 $X=8456000 $Y=9376000
X3473 3436 24 aoi22 $T=8464000 2880000 0 0 $X=8464000 $Y=2880000
X3474 3437 24 aoi22 $T=8472000 9608000 0 0 $X=8472000 $Y=9608000
X3475 3438 24 aoi22 $T=8480000 6360000 0 0 $X=8480000 $Y=6360000
X3476 3439 24 aoi22 $T=8512000 4504000 0 0 $X=8512000 $Y=4504000
X3477 3440 24 aoi22 $T=8520000 13088000 0 0 $X=8520000 $Y=13088000
X3478 3441 24 aoi22 $T=8536000 328000 0 0 $X=8536000 $Y=328000
X3479 3442 24 aoi22 $T=8536000 4968000 0 0 $X=8536000 $Y=4968000
X3480 3443 24 aoi22 $T=8536000 6360000 0 0 $X=8536000 $Y=6360000
X3481 3444 24 aoi22 $T=8608000 9840000 0 0 $X=8608000 $Y=9840000
X3482 3445 24 aoi22 $T=8656000 4968000 0 0 $X=8656000 $Y=4968000
X3483 3446 24 aoi22 $T=8688000 8680000 0 0 $X=8688000 $Y=8680000
X3484 3447 24 aoi22 $T=8745000 11000000 1 180 $X=8696000 $Y=11000000
X3485 3448 24 aoi22 $T=8744000 7752000 0 0 $X=8744000 $Y=7752000
X3486 3449 24 aoi22 $T=8752000 13320000 0 0 $X=8752000 $Y=13320000
X3487 3450 24 aoi22 $T=8760000 9376000 0 0 $X=8760000 $Y=9376000
X3488 3451 24 aoi22 $T=8776000 7056000 0 0 $X=8776000 $Y=7056000
X3489 3452 24 aoi22 $T=8841000 3576000 1 180 $X=8792000 $Y=3576000
X3490 3453 24 aoi22 $T=8792000 7520000 0 0 $X=8792000 $Y=7520000
X3491 3454 24 aoi22 $T=8857000 8216000 1 180 $X=8808000 $Y=8216000
X3492 3455 24 aoi22 $T=8808000 13320000 0 0 $X=8808000 $Y=13320000
X3493 3456 24 aoi22 $T=8816000 8448000 0 0 $X=8816000 $Y=8448000
X3494 3457 24 aoi22 $T=8824000 13088000 0 0 $X=8824000 $Y=13088000
X3495 3458 24 aoi22 $T=8881000 11696000 1 180 $X=8832000 $Y=11696000
X3496 3459 24 aoi22 $T=8840000 4736000 0 0 $X=8840000 $Y=4736000
X3497 3460 24 aoi22 $T=8864000 13320000 0 0 $X=8864000 $Y=13320000
X3498 3461 24 aoi22 $T=8945000 3344000 1 180 $X=8896000 $Y=3344000
X3499 3462 24 aoi22 $T=8993000 11696000 1 180 $X=8944000 $Y=11696000
X3500 3463 24 aoi22 $T=8992000 1256000 0 0 $X=8992000 $Y=1256000
X3501 3464 24 aoi22 $T=9016000 11464000 0 0 $X=9016000 $Y=11464000
X3502 3465 24 aoi22 $T=9065000 12392000 1 180 $X=9016000 $Y=12392000
X3503 3466 24 aoi22 $T=9113000 4504000 1 180 $X=9064000 $Y=4504000
X3504 3467 24 aoi22 $T=9113000 8912000 1 180 $X=9064000 $Y=8912000
X3505 3468 24 aoi22 $T=9113000 9840000 1 180 $X=9064000 $Y=9840000
X3506 3469 24 aoi22 $T=9064000 12160000 0 0 $X=9064000 $Y=12160000
X3507 3470 24 aoi22 $T=9104000 4272000 0 0 $X=9104000 $Y=4272000
X3508 3471 24 aoi22 $T=9161000 7056000 1 180 $X=9112000 $Y=7056000
X3509 3472 24 aoi22 $T=9112000 11928000 0 0 $X=9112000 $Y=11928000
X3510 3473 24 aoi22 $T=9120000 1024000 0 0 $X=9120000 $Y=1024000
X3511 3474 24 aoi22 $T=9120000 12160000 0 0 $X=9120000 $Y=12160000
X3512 3475 24 aoi22 $T=9128000 10304000 0 0 $X=9128000 $Y=10304000
X3513 3476 24 aoi22 $T=9128000 12392000 0 0 $X=9128000 $Y=12392000
X3514 3477 24 aoi22 $T=9152000 10536000 0 0 $X=9152000 $Y=10536000
X3515 3478 24 aoi22 $T=9176000 1024000 0 0 $X=9176000 $Y=1024000
X3516 3479 24 aoi22 $T=9176000 8912000 0 0 $X=9176000 $Y=8912000
X3517 3480 24 aoi22 $T=9200000 6360000 0 0 $X=9200000 $Y=6360000
X3518 3481 24 aoi22 $T=9208000 4736000 0 0 $X=9208000 $Y=4736000
X3519 3482 24 aoi22 $T=9289000 7984000 1 180 $X=9240000 $Y=7984000
X3520 3483 24 aoi22 $T=9313000 7288000 1 180 $X=9264000 $Y=7288000
X3521 3484 24 aoi22 $T=9272000 9840000 0 0 $X=9272000 $Y=9840000
X3522 3485 24 aoi22 $T=9280000 7520000 0 0 $X=9280000 $Y=7520000
X3523 3486 24 aoi22 $T=9296000 4040000 0 0 $X=9296000 $Y=4040000
X3524 3487 24 aoi22 $T=9296000 5664000 0 0 $X=9296000 $Y=5664000
X3525 3488 24 aoi22 $T=9401000 4040000 1 180 $X=9352000 $Y=4040000
X3526 3489 24 aoi22 $T=9360000 1256000 0 0 $X=9360000 $Y=1256000
X3527 3490 24 aoi22 $T=9409000 7984000 1 180 $X=9360000 $Y=7984000
X3528 3491 24 aoi22 $T=9456000 1952000 0 0 $X=9456000 $Y=1952000
X3529 3492 24 aoi22 $T=9464000 4040000 0 0 $X=9464000 $Y=4040000
X3530 3493 24 aoi22 $T=9480000 1256000 0 0 $X=9480000 $Y=1256000
X3531 3494 24 aoi22 $T=9496000 9376000 0 0 $X=9496000 $Y=9376000
X3532 3495 24 aoi22 $T=9504000 3808000 0 0 $X=9504000 $Y=3808000
X3533 3496 24 aoi22 $T=9512000 1952000 0 0 $X=9512000 $Y=1952000
X3534 3497 24 aoi22 $T=9520000 4040000 0 0 $X=9520000 $Y=4040000
X3535 3498 24 aoi22 $T=9536000 792000 0 0 $X=9536000 $Y=792000
X3536 3499 24 aoi22 $T=9585000 8912000 1 180 $X=9536000 $Y=8912000
X3537 3500 24 aoi22 $T=9576000 4040000 0 0 $X=9576000 $Y=4040000
X3538 3501 24 aoi22 $T=9600000 560000 0 0 $X=9600000 $Y=560000
X3539 3502 24 aoi22 $T=9681000 4040000 1 180 $X=9632000 $Y=4040000
X3540 3503 24 aoi22 $T=9713000 7984000 1 180 $X=9664000 $Y=7984000
X3541 3504 24 aoi22 $T=9745000 1720000 1 180 $X=9696000 $Y=1720000
X3542 3505 24 aoi22 $T=9753000 10536000 1 180 $X=9704000 $Y=10536000
X3543 3506 24 aoi22 $T=9769000 8216000 1 180 $X=9720000 $Y=8216000
X3544 3507 24 aoi22 $T=9785000 9608000 1 180 $X=9736000 $Y=9608000
X3545 3508 24 aoi22 $T=9752000 328000 0 0 $X=9752000 $Y=328000
X3546 3509 24 aoi22 $T=9801000 10768000 1 180 $X=9752000 $Y=10768000
X3547 3510 24 aoi22 $T=9760000 2648000 0 0 $X=9760000 $Y=2648000
X3548 3511 24 aoi22 $T=9768000 6592000 0 0 $X=9768000 $Y=6592000
X3549 3512 24 aoi22 $T=9776000 8216000 0 0 $X=9776000 $Y=8216000
X3550 3513 24 aoi22 $T=9849000 11696000 1 180 $X=9800000 $Y=11696000
X3551 3514 24 aoi22 $T=9808000 8680000 0 0 $X=9808000 $Y=8680000
X3552 3515 24 aoi22 $T=9824000 2184000 0 0 $X=9824000 $Y=2184000
X3553 3516 24 aoi22 $T=9929000 7056000 1 180 $X=9880000 $Y=7056000
X3554 3517 24 aoi22 $T=9937000 5896000 1 180 $X=9888000 $Y=5896000
X3555 3518 24 aoi22 $T=9945000 4504000 1 180 $X=9896000 $Y=4504000
X3556 3519 24 aoi22 $T=9904000 10768000 0 0 $X=9904000 $Y=10768000
X3557 3520 24 aoi22 $T=9993000 5896000 1 180 $X=9944000 $Y=5896000
X3558 3521 24 aoi22 $T=10025000 1024000 1 180 $X=9976000 $Y=1024000
X3559 3522 24 aoi22 $T=9992000 4040000 0 0 $X=9992000 $Y=4040000
X3560 3523 24 aoi22 $T=10000000 5896000 0 0 $X=10000000 $Y=5896000
X3561 3524 24 aoi22 $T=10000000 10536000 0 0 $X=10000000 $Y=10536000
X3562 3525 24 aoi22 $T=10057000 9144000 1 180 $X=10008000 $Y=9144000
X3563 3526 24 aoi22 $T=10024000 7984000 0 0 $X=10024000 $Y=7984000
X3564 3527 24 aoi22 $T=10040000 9608000 0 0 $X=10040000 $Y=9608000
X3565 3528 24 aoi22 $T=10048000 4040000 0 0 $X=10048000 $Y=4040000
X3566 3529 24 aoi22 $T=10105000 6360000 1 180 $X=10056000 $Y=6360000
X3567 3530 24 aoi22 $T=10113000 9144000 1 180 $X=10064000 $Y=9144000
X3568 3531 24 aoi22 $T=10088000 1024000 0 0 $X=10088000 $Y=1024000
X3569 3532 24 aoi22 $T=10137000 13320000 1 180 $X=10088000 $Y=13320000
X3570 3533 24 aoi22 $T=10152000 5200000 0 0 $X=10152000 $Y=5200000
X3571 3534 24 aoi22 $T=10208000 9144000 0 0 $X=10208000 $Y=9144000
X3572 2352 24 aoi22 $T=10265000 5664000 1 180 $X=10216000 $Y=5664000
X3573 3535 24 aoi22 $T=10240000 11000000 0 0 $X=10240000 $Y=11000000
X3574 3536 24 aoi22 $T=10248000 11928000 0 0 $X=10248000 $Y=11928000
X3575 3537 24 aoi22 $T=10305000 4504000 1 180 $X=10256000 $Y=4504000
X3576 3538 24 aoi22 $T=10264000 9144000 0 0 $X=10264000 $Y=9144000
X3577 3539 24 aoi22 $T=10313000 12392000 1 180 $X=10264000 $Y=12392000
X3578 3540 24 aoi22 $T=10264000 13320000 0 0 $X=10264000 $Y=13320000
X3579 3541 24 aoi22 $T=10337000 3112000 1 180 $X=10288000 $Y=3112000
X3580 3542 24 aoi22 $T=10353000 1952000 1 180 $X=10304000 $Y=1952000
X3581 3543 24 aoi22 $T=10353000 10536000 1 180 $X=10304000 $Y=10536000
X3582 3544 24 aoi22 $T=10320000 9144000 0 0 $X=10320000 $Y=9144000
X3583 3545 24 aoi22 $T=10336000 5664000 0 0 $X=10336000 $Y=5664000
X3584 3546 24 aoi22 $T=10368000 2648000 0 0 $X=10368000 $Y=2648000
X3585 3547 24 aoi22 $T=10376000 2184000 0 0 $X=10376000 $Y=2184000
X3586 3548 24 aoi22 $T=10376000 6592000 0 0 $X=10376000 $Y=6592000
X3587 3549 24 aoi22 $T=10376000 9144000 0 0 $X=10376000 $Y=9144000
X3588 3550 24 aoi22 $T=10376000 12392000 0 0 $X=10376000 $Y=12392000
X3589 3551 24 aoi22 $T=10416000 1952000 0 0 $X=10416000 $Y=1952000
X3590 3552 24 aoi22 $T=10424000 2648000 0 0 $X=10424000 $Y=2648000
X3591 3553 24 aoi22 $T=10432000 2880000 0 0 $X=10432000 $Y=2880000
X3592 3554 24 aoi22 $T=10464000 560000 0 0 $X=10464000 $Y=560000
X3593 3555 24 aoi22 $T=10513000 2184000 1 180 $X=10464000 $Y=2184000
X3594 3556 24 aoi22 $T=10521000 8912000 1 180 $X=10472000 $Y=8912000
X3595 3557 24 aoi22 $T=10488000 11464000 0 0 $X=10488000 $Y=11464000
X3596 3558 24 aoi22 $T=10520000 3344000 0 0 $X=10520000 $Y=3344000
X3597 3559 24 aoi22 $T=10528000 8912000 0 0 $X=10528000 $Y=8912000
X3598 3560 24 aoi22 $T=10544000 7056000 0 0 $X=10544000 $Y=7056000
X3599 3561 24 aoi22 $T=10544000 11464000 0 0 $X=10544000 $Y=11464000
X3600 3562 24 aoi22 $T=10584000 3576000 0 0 $X=10584000 $Y=3576000
X3601 3563 24 aoi22 $T=10640000 8912000 0 0 $X=10640000 $Y=8912000
X3602 3564 24 aoi22 $T=10640000 11696000 0 0 $X=10640000 $Y=11696000
X3603 3565 24 aoi22 $T=10672000 10536000 0 0 $X=10672000 $Y=10536000
X3604 3566 24 aoi22 $T=10688000 4736000 0 0 $X=10688000 $Y=4736000
X3605 3567 24 aoi22 $T=10704000 3576000 0 0 $X=10704000 $Y=3576000
X3606 3568 24 aoi22 $T=10712000 9840000 0 0 $X=10712000 $Y=9840000
X3607 3569 24 aoi22 $T=10769000 4504000 1 180 $X=10720000 $Y=4504000
X3608 3570 24 aoi22 $T=10728000 10536000 0 0 $X=10728000 $Y=10536000
X3609 3571 24 aoi22 $T=10736000 9608000 0 0 $X=10736000 $Y=9608000
X3610 3572 24 aoi22 $T=10744000 6128000 0 0 $X=10744000 $Y=6128000
X3611 3573 24 aoi22 $T=10825000 6824000 1 180 $X=10776000 $Y=6824000
X3612 3574 24 aoi22 $T=10776000 13320000 0 0 $X=10776000 $Y=13320000
X3613 3575 24 aoi22 $T=10792000 7984000 0 0 $X=10792000 $Y=7984000
X3614 3576 24 aoi22 $T=10792000 12856000 0 0 $X=10792000 $Y=12856000
X3615 3577 24 aoi22 $T=10849000 10768000 1 180 $X=10800000 $Y=10768000
X3616 3578 24 aoi22 $T=10857000 7752000 1 180 $X=10808000 $Y=7752000
X3617 3579 24 aoi22 $T=10808000 8216000 0 0 $X=10808000 $Y=8216000
X3618 3580 24 aoi22 $T=10808000 9376000 0 0 $X=10808000 $Y=9376000
X3619 3581 24 aoi22 $T=10808000 11696000 0 0 $X=10808000 $Y=11696000
X3620 3582 24 aoi22 $T=10865000 5200000 1 180 $X=10816000 $Y=5200000
X3621 3583 24 aoi22 $T=10832000 4504000 0 0 $X=10832000 $Y=4504000
X3622 3584 24 aoi22 $T=10840000 13088000 0 0 $X=10840000 $Y=13088000
X3623 3585 24 aoi22 $T=10856000 5896000 0 0 $X=10856000 $Y=5896000
X3624 3586 24 aoi22 $T=10856000 6128000 0 0 $X=10856000 $Y=6128000
X3625 3587 24 aoi22 $T=10864000 9376000 0 0 $X=10864000 $Y=9376000
X3626 3588 24 aoi22 $T=10880000 2184000 0 0 $X=10880000 $Y=2184000
X3627 3589 24 aoi22 $T=10880000 5664000 0 0 $X=10880000 $Y=5664000
X3628 3590 24 aoi22 $T=10888000 11000000 0 0 $X=10888000 $Y=11000000
X3629 3591 24 aoi22 $T=10904000 792000 0 0 $X=10904000 $Y=792000
X3630 3592 24 aoi22 $T=10920000 8216000 0 0 $X=10920000 $Y=8216000
X3631 3593 24 aoi22 $T=10936000 2184000 0 0 $X=10936000 $Y=2184000
X3632 3594 24 aoi22 $T=10976000 8216000 0 0 $X=10976000 $Y=8216000
X3633 3595 24 aoi22 $T=10992000 13088000 0 0 $X=10992000 $Y=13088000
X3634 3596 24 aoi22 $T=10992000 13320000 0 0 $X=10992000 $Y=13320000
X3635 3597 24 aoi22 $T=11032000 8216000 0 0 $X=11032000 $Y=8216000
X3636 3598 24 aoi22 $T=11048000 11232000 0 0 $X=11048000 $Y=11232000
X3637 3599 24 aoi22 $T=11072000 3576000 0 0 $X=11072000 $Y=3576000
X3638 3600 24 aoi22 $T=11088000 10536000 0 0 $X=11088000 $Y=10536000
X3639 3601 24 aoi22 $T=11120000 5432000 0 0 $X=11120000 $Y=5432000
X3640 3602 24 aoi22 $T=11144000 10536000 0 0 $X=11144000 $Y=10536000
X3641 3603 24 aoi22 $T=11289000 9144000 1 180 $X=11240000 $Y=9144000
X3642 3604 24 aoi22 $T=11256000 10536000 0 0 $X=11256000 $Y=10536000
X3643 3605 24 aoi22 $T=11321000 3808000 1 180 $X=11272000 $Y=3808000
X3644 3606 24 aoi22 $T=11321000 4736000 1 180 $X=11272000 $Y=4736000
X3645 3607 24 aoi22 $T=11288000 9608000 0 0 $X=11288000 $Y=9608000
X3646 3608 24 aoi22 $T=11312000 10536000 0 0 $X=11312000 $Y=10536000
X3647 3609 24 aoi22 $T=11377000 4736000 1 180 $X=11328000 $Y=4736000
X3648 3610 24 aoi22 $T=11328000 9840000 0 0 $X=11328000 $Y=9840000
X3649 3611 24 aoi22 $T=11344000 5896000 0 0 $X=11344000 $Y=5896000
X3650 3612 24 aoi22 $T=11409000 7752000 1 180 $X=11360000 $Y=7752000
X3651 3613 24 aoi22 $T=11368000 10536000 0 0 $X=11368000 $Y=10536000
X3652 3614 24 aoi22 $T=11425000 3576000 1 180 $X=11376000 $Y=3576000
X3653 3615 24 aoi22 $T=11425000 7984000 1 180 $X=11376000 $Y=7984000
X3654 3616 24 aoi22 $T=11384000 9840000 0 0 $X=11384000 $Y=9840000
X3655 3617 24 aoi22 $T=11416000 9608000 0 0 $X=11416000 $Y=9608000
X3656 3618 24 aoi22 $T=11424000 5200000 0 0 $X=11424000 $Y=5200000
X3657 3619 24 aoi22 $T=11424000 10536000 0 0 $X=11424000 $Y=10536000
X3658 3620 24 aoi22 $T=11432000 12624000 0 0 $X=11432000 $Y=12624000
X3659 3621 24 aoi22 $T=11440000 4736000 0 0 $X=11440000 $Y=4736000
X3660 3622 24 aoi22 $T=11472000 7752000 0 0 $X=11472000 $Y=7752000
X3661 3623 24 aoi22 $T=11472000 9608000 0 0 $X=11472000 $Y=9608000
X3662 3624 24 aoi22 $T=11480000 5200000 0 0 $X=11480000 $Y=5200000
X3663 3625 24 aoi22 $T=11480000 5432000 0 0 $X=11480000 $Y=5432000
X3664 3626 24 aoi22 $T=11537000 2416000 1 180 $X=11488000 $Y=2416000
X3665 3627 24 aoi22 $T=11496000 3344000 0 0 $X=11496000 $Y=3344000
X3666 3628 24 aoi22 $T=11545000 7984000 1 180 $X=11496000 $Y=7984000
X3667 3629 24 aoi22 $T=11496000 10072000 0 0 $X=11496000 $Y=10072000
X3668 3630 24 aoi22 $T=11520000 12392000 0 0 $X=11520000 $Y=12392000
X3669 3631 24 aoi22 $T=11577000 7752000 1 180 $X=11528000 $Y=7752000
X3670 3632 24 aoi22 $T=11577000 11696000 1 180 $X=11528000 $Y=11696000
X3671 3633 24 aoi22 $T=11544000 12624000 0 0 $X=11544000 $Y=12624000
X3672 3634 24 aoi22 $T=11552000 11000000 0 0 $X=11552000 $Y=11000000
X3673 3635 24 aoi22 $T=11568000 3808000 0 0 $X=11568000 $Y=3808000
X3674 3636 24 aoi22 $T=11600000 10768000 0 0 $X=11600000 $Y=10768000
X3675 3637 24 aoi22 $T=11600000 12624000 0 0 $X=11600000 $Y=12624000
X3676 3638 24 aoi22 $T=11608000 6360000 0 0 $X=11608000 $Y=6360000
X3677 3639 24 aoi22 $T=11608000 11000000 0 0 $X=11608000 $Y=11000000
X3678 3640 24 aoi22 $T=11616000 1952000 0 0 $X=11616000 $Y=1952000
X3679 3641 24 aoi22 $T=11665000 6824000 1 180 $X=11616000 $Y=6824000
X3680 3642 24 aoi22 $T=11624000 2648000 0 0 $X=11624000 $Y=2648000
X3681 3643 24 aoi22 $T=11624000 3808000 0 0 $X=11624000 $Y=3808000
X3682 3644 24 aoi22 $T=11632000 12392000 0 0 $X=11632000 $Y=12392000
X3683 3645 24 aoi22 $T=11640000 7752000 0 0 $X=11640000 $Y=7752000
X3684 3646 24 aoi22 $T=11640000 11696000 0 0 $X=11640000 $Y=11696000
X3685 3647 24 aoi22 $T=11656000 12624000 0 0 $X=11656000 $Y=12624000
X3686 3648 24 aoi22 $T=11664000 11232000 0 0 $X=11664000 $Y=11232000
X3687 3649 24 aoi22 $T=11672000 1952000 0 0 $X=11672000 $Y=1952000
X3688 3650 24 aoi22 $T=11688000 6592000 0 0 $X=11688000 $Y=6592000
X3689 3651 24 aoi22 $T=11712000 12624000 0 0 $X=11712000 $Y=12624000
X3690 3652 24 aoi22 $T=11728000 4040000 0 0 $X=11728000 $Y=4040000
X3691 3653 24 aoi22 $T=11792000 7752000 0 0 $X=11792000 $Y=7752000
X3692 3654 24 aoi22 $T=11800000 6592000 0 0 $X=11800000 $Y=6592000
X3693 3655 24 aoi22 $T=11856000 6592000 0 0 $X=11856000 $Y=6592000
X3694 3656 24 aoi22 $T=11912000 6592000 0 0 $X=11912000 $Y=6592000
X3695 3657 24 aoi22 $T=11976000 2184000 0 0 $X=11976000 $Y=2184000
X3696 3658 24 aoi22 $T=12033000 3112000 1 180 $X=11984000 $Y=3112000
X3697 3659 24 aoi22 $T=12040000 3112000 0 0 $X=12040000 $Y=3112000
X3698 3660 24 aoi22 $T=12040000 11464000 0 0 $X=12040000 $Y=11464000
X3699 3661 24 aoi22 $T=12104000 3576000 0 0 $X=12104000 $Y=3576000
X3700 3662 24 aoi22 $T=12168000 3808000 0 0 $X=12168000 $Y=3808000
X3701 3663 24 aoi22 $T=12224000 3808000 0 0 $X=12224000 $Y=3808000
X3702 3664 24 aoi22 $T=12224000 4736000 0 0 $X=12224000 $Y=4736000
X3703 24 3665 ICV_1 $T=336000 5432000 1 180 $X=152000 $Y=5432000
X3704 24 3666 ICV_1 $T=336000 9144000 1 180 $X=152000 $Y=9144000
X3705 24 3667 ICV_1 $T=336000 9376000 1 180 $X=152000 $Y=9376000
X3706 24 3668 ICV_1 $T=336000 11000000 1 180 $X=152000 $Y=11000000
X3707 24 3669 ICV_1 $T=376000 7752000 1 180 $X=192000 $Y=7752000
X3708 24 3670 ICV_1 $T=584000 6824000 1 180 $X=400000 $Y=6824000
X3709 24 3671 ICV_1 $T=640000 6128000 1 180 $X=456000 $Y=6128000
X3710 24 3672 ICV_1 $T=704000 5432000 1 180 $X=520000 $Y=5432000
X3711 24 3673 ICV_1 $T=824000 12392000 1 180 $X=640000 $Y=12392000
X3712 24 3674 ICV_1 $T=832000 6824000 1 180 $X=648000 $Y=6824000
X3713 24 3675 ICV_1 $T=872000 12856000 1 180 $X=688000 $Y=12856000
X3714 24 3676 ICV_1 $T=888000 7288000 1 180 $X=704000 $Y=7288000
X3715 24 3677 ICV_1 $T=1064000 6128000 1 180 $X=880000 $Y=6128000
X3716 24 3678 ICV_1 $T=1064000 9376000 1 180 $X=880000 $Y=9376000
X3717 24 3679 ICV_1 $T=1136000 5200000 1 180 $X=952000 $Y=5200000
X3718 24 3680 ICV_1 $T=1144000 6824000 1 180 $X=960000 $Y=6824000
X3719 24 3681 ICV_1 $T=1160000 8216000 1 180 $X=976000 $Y=8216000
X3720 24 3682 ICV_1 $T=1256000 5896000 1 180 $X=1072000 $Y=5896000
X3721 24 3683 ICV_1 $T=1272000 4272000 1 180 $X=1088000 $Y=4272000
X3722 24 3684 ICV_1 $T=1304000 7056000 1 180 $X=1120000 $Y=7056000
X3723 24 3685 ICV_1 $T=1352000 7288000 1 180 $X=1168000 $Y=7288000
X3724 24 3686 ICV_1 $T=1392000 6824000 1 180 $X=1208000 $Y=6824000
X3725 24 3687 ICV_1 $T=1392000 13552000 1 180 $X=1208000 $Y=13552000
X3726 24 3688 ICV_1 $T=1408000 7520000 1 180 $X=1224000 $Y=7520000
X3727 24 3689 ICV_1 $T=1440000 4504000 1 180 $X=1256000 $Y=4504000
X3728 24 3690 ICV_1 $T=1440000 6360000 1 180 $X=1256000 $Y=6360000
X3729 24 3691 ICV_1 $T=1440000 8216000 1 180 $X=1256000 $Y=8216000
X3730 24 3692 ICV_1 $T=1448000 4736000 1 180 $X=1264000 $Y=4736000
X3731 24 3693 ICV_1 $T=1448000 8448000 1 180 $X=1264000 $Y=8448000
X3732 24 3694 ICV_1 $T=1456000 7752000 1 180 $X=1272000 $Y=7752000
X3733 24 3695 ICV_1 $T=1464000 4968000 1 180 $X=1280000 $Y=4968000
X3734 24 3696 ICV_1 $T=1464000 9376000 1 180 $X=1280000 $Y=9376000
X3735 24 3697 ICV_1 $T=1472000 6128000 1 180 $X=1288000 $Y=6128000
X3736 24 3698 ICV_1 $T=1496000 7984000 1 180 $X=1312000 $Y=7984000
X3737 24 3699 ICV_1 $T=1512000 5432000 1 180 $X=1328000 $Y=5432000
X3738 24 3700 ICV_1 $T=1520000 4272000 1 180 $X=1336000 $Y=4272000
X3739 24 3701 ICV_1 $T=1536000 5896000 1 180 $X=1352000 $Y=5896000
X3740 24 3702 ICV_1 $T=1536000 8912000 1 180 $X=1352000 $Y=8912000
X3741 24 3703 ICV_1 $T=1544000 8680000 1 180 $X=1360000 $Y=8680000
X3742 24 3704 ICV_1 $T=1552000 9144000 1 180 $X=1368000 $Y=9144000
X3743 24 3705 ICV_1 $T=1592000 5664000 1 180 $X=1408000 $Y=5664000
X3744 24 3706 ICV_1 $T=1696000 4504000 1 180 $X=1512000 $Y=4504000
X3745 24 3707 ICV_1 $T=1696000 9608000 1 180 $X=1512000 $Y=9608000
X3746 24 3708 ICV_1 $T=1728000 4736000 1 180 $X=1544000 $Y=4736000
X3747 24 3709 ICV_1 $T=1768000 4272000 1 180 $X=1584000 $Y=4272000
X3748 24 3710 ICV_1 $T=1856000 12624000 1 180 $X=1672000 $Y=12624000
X3749 24 3711 ICV_1 $T=1984000 11000000 1 180 $X=1800000 $Y=11000000
X3750 24 3712 ICV_1 $T=2016000 12160000 1 180 $X=1832000 $Y=12160000
X3751 24 3713 ICV_1 $T=2024000 9376000 1 180 $X=1840000 $Y=9376000
X3752 24 3714 ICV_1 $T=2032000 11464000 1 180 $X=1848000 $Y=11464000
X3753 24 3715 ICV_1 $T=2056000 7984000 1 180 $X=1872000 $Y=7984000
X3754 24 3716 ICV_1 $T=2072000 12856000 1 180 $X=1888000 $Y=12856000
X3755 24 3717 ICV_1 $T=2088000 4736000 1 180 $X=1904000 $Y=4736000
X3756 24 3718 ICV_1 $T=2104000 10768000 1 180 $X=1920000 $Y=10768000
X3757 24 3719 ICV_1 $T=2152000 7056000 1 180 $X=1968000 $Y=7056000
X3758 24 3720 ICV_1 $T=2160000 7752000 1 180 $X=1976000 $Y=7752000
X3759 24 3721 ICV_1 $T=2248000 5432000 1 180 $X=2064000 $Y=5432000
X3760 24 3722 ICV_1 $T=2280000 12392000 1 180 $X=2096000 $Y=12392000
X3761 24 3723 ICV_1 $T=2288000 9840000 1 180 $X=2104000 $Y=9840000
X3762 24 3724 ICV_1 $T=2320000 11232000 1 180 $X=2136000 $Y=11232000
X3763 24 3725 ICV_1 $T=2344000 4040000 1 180 $X=2160000 $Y=4040000
X3764 24 3726 ICV_1 $T=2392000 10768000 1 180 $X=2208000 $Y=10768000
X3765 24 3727 ICV_1 $T=2424000 12160000 1 180 $X=2240000 $Y=12160000
X3766 24 3728 ICV_1 $T=2496000 8912000 1 180 $X=2312000 $Y=8912000
X3767 24 3729 ICV_1 $T=2600000 13088000 1 180 $X=2416000 $Y=13088000
X3768 24 3730 ICV_1 $T=2608000 9376000 1 180 $X=2424000 $Y=9376000
X3769 24 3731 ICV_1 $T=2608000 9840000 1 180 $X=2424000 $Y=9840000
X3770 24 3732 ICV_1 $T=2672000 3576000 1 180 $X=2488000 $Y=3576000
X3771 24 3733 ICV_1 $T=2672000 11464000 1 180 $X=2488000 $Y=11464000
X3772 24 3734 ICV_1 $T=2696000 10072000 1 180 $X=2512000 $Y=10072000
X3773 24 3735 ICV_1 $T=2728000 3808000 1 180 $X=2544000 $Y=3808000
X3774 24 3736 ICV_1 $T=2760000 11232000 1 180 $X=2576000 $Y=11232000
X3775 24 3737 ICV_1 $T=2768000 10768000 1 180 $X=2584000 $Y=10768000
X3776 24 3738 ICV_1 $T=2800000 4968000 1 180 $X=2616000 $Y=4968000
X3777 24 3739 ICV_1 $T=2832000 6592000 1 180 $X=2648000 $Y=6592000
X3778 24 3740 ICV_1 $T=2848000 7984000 1 180 $X=2664000 $Y=7984000
X3779 24 3741 ICV_1 $T=2856000 9840000 1 180 $X=2672000 $Y=9840000
X3780 24 3742 ICV_1 $T=2904000 9608000 1 180 $X=2720000 $Y=9608000
X3781 24 3743 ICV_1 $T=2920000 12624000 1 180 $X=2736000 $Y=12624000
X3782 24 3744 ICV_1 $T=2928000 6128000 1 180 $X=2744000 $Y=6128000
X3783 24 3745 ICV_1 $T=2936000 3112000 1 180 $X=2752000 $Y=3112000
X3784 24 3746 ICV_1 $T=2968000 6360000 1 180 $X=2784000 $Y=6360000
X3785 24 3747 ICV_1 $T=2984000 9376000 1 180 $X=2800000 $Y=9376000
X3786 24 3748 ICV_1 $T=3008000 7520000 1 180 $X=2824000 $Y=7520000
X3787 24 3749 ICV_1 $T=3112000 8912000 1 180 $X=2928000 $Y=8912000
X3788 24 3750 ICV_1 $T=3120000 8448000 1 180 $X=2936000 $Y=8448000
X3789 24 3751 ICV_1 $T=3152000 9608000 1 180 $X=2968000 $Y=9608000
X3790 24 3752 ICV_1 $T=3160000 8680000 1 180 $X=2976000 $Y=8680000
X3791 24 3753 ICV_1 $T=3184000 5896000 1 180 $X=3000000 $Y=5896000
X3792 24 3754 ICV_1 $T=3200000 11464000 1 180 $X=3016000 $Y=11464000
X3793 24 3755 ICV_1 $T=3208000 9144000 1 180 $X=3024000 $Y=9144000
X3794 24 3756 ICV_1 $T=3352000 3808000 1 180 $X=3168000 $Y=3808000
X3795 24 3757 ICV_1 $T=3376000 11928000 1 180 $X=3192000 $Y=11928000
X3796 24 3758 ICV_1 $T=3408000 8680000 1 180 $X=3224000 $Y=8680000
X3797 24 3759 ICV_1 $T=3560000 11000000 1 180 $X=3376000 $Y=11000000
X3798 24 3760 ICV_1 $T=3608000 11232000 1 180 $X=3424000 $Y=11232000
X3799 24 3761 ICV_1 $T=3608000 13088000 1 180 $X=3424000 $Y=13088000
X3800 24 3762 ICV_1 $T=3616000 8216000 1 180 $X=3432000 $Y=8216000
X3801 24 3763 ICV_1 $T=3616000 13552000 1 180 $X=3432000 $Y=13552000
X3802 24 3764 ICV_1 $T=3648000 8448000 1 180 $X=3464000 $Y=8448000
X3803 24 3765 ICV_1 $T=3664000 6592000 1 180 $X=3480000 $Y=6592000
X3804 24 3766 ICV_1 $T=3680000 12392000 1 180 $X=3496000 $Y=12392000
X3805 24 3767 ICV_1 $T=3688000 13320000 1 180 $X=3504000 $Y=13320000
X3806 24 3768 ICV_1 $T=3760000 11464000 1 180 $X=3576000 $Y=11464000
X3807 24 3769 ICV_1 $T=3808000 9840000 1 180 $X=3624000 $Y=9840000
X3808 24 3770 ICV_1 $T=3816000 9608000 1 180 $X=3632000 $Y=9608000
X3809 24 3771 ICV_1 $T=3912000 11232000 1 180 $X=3728000 $Y=11232000
X3810 24 3772 ICV_1 $T=3928000 10072000 1 180 $X=3744000 $Y=10072000
X3811 24 3773 ICV_1 $T=3944000 7984000 1 180 $X=3760000 $Y=7984000
X3812 24 3774 ICV_1 $T=3976000 5664000 1 180 $X=3792000 $Y=5664000
X3813 24 3775 ICV_1 $T=3976000 6360000 1 180 $X=3792000 $Y=6360000
X3814 24 3776 ICV_1 $T=4000000 6128000 1 180 $X=3816000 $Y=6128000
X3815 24 3777 ICV_1 $T=4040000 5896000 1 180 $X=3856000 $Y=5896000
X3816 24 3778 ICV_1 $T=4088000 4504000 1 180 $X=3904000 $Y=4504000
X3817 24 3779 ICV_1 $T=4192000 7984000 1 180 $X=4008000 $Y=7984000
X3818 24 3780 ICV_1 $T=4216000 9608000 1 180 $X=4032000 $Y=9608000
X3819 24 3781 ICV_1 $T=4240000 2184000 1 180 $X=4056000 $Y=2184000
X3820 24 3782 ICV_1 $T=4248000 10072000 1 180 $X=4064000 $Y=10072000
X3821 24 3783 ICV_1 $T=4280000 4040000 1 180 $X=4096000 $Y=4040000
X3822 24 3784 ICV_1 $T=4288000 7288000 1 180 $X=4104000 $Y=7288000
X3823 24 3785 ICV_1 $T=4288000 13088000 1 180 $X=4104000 $Y=13088000
X3824 24 3786 ICV_1 $T=4296000 12160000 1 180 $X=4112000 $Y=12160000
X3825 24 3787 ICV_1 $T=4296000 12392000 1 180 $X=4112000 $Y=12392000
X3826 24 3788 ICV_1 $T=4328000 12856000 1 180 $X=4144000 $Y=12856000
X3827 24 3789 ICV_1 $T=4336000 11928000 1 180 $X=4152000 $Y=11928000
X3828 24 3790 ICV_1 $T=4344000 7056000 1 180 $X=4160000 $Y=7056000
X3829 24 3791 ICV_1 $T=4344000 11696000 1 180 $X=4160000 $Y=11696000
X3830 24 3792 ICV_1 $T=4368000 6824000 1 180 $X=4184000 $Y=6824000
X3831 24 3793 ICV_1 $T=4424000 3112000 1 180 $X=4240000 $Y=3112000
X3832 24 3794 ICV_1 $T=4464000 13552000 1 180 $X=4280000 $Y=13552000
X3833 24 3795 ICV_1 $T=4480000 560000 1 180 $X=4296000 $Y=560000
X3834 24 3796 ICV_1 $T=4496000 10072000 1 180 $X=4312000 $Y=10072000
X3835 24 3797 ICV_1 $T=4520000 6592000 1 180 $X=4336000 $Y=6592000
X3836 24 3798 ICV_1 $T=4520000 7752000 1 180 $X=4336000 $Y=7752000
X3837 24 3799 ICV_1 $T=4528000 7984000 1 180 $X=4344000 $Y=7984000
X3838 24 3800 ICV_1 $T=4536000 792000 1 180 $X=4352000 $Y=792000
X3839 24 3801 ICV_1 $T=4568000 9376000 1 180 $X=4384000 $Y=9376000
X3840 24 3802 ICV_1 $T=4576000 8912000 1 180 $X=4392000 $Y=8912000
X3841 24 3803 ICV_1 $T=4584000 4968000 1 180 $X=4400000 $Y=4968000
X3842 24 3804 ICV_1 $T=4592000 7056000 1 180 $X=4408000 $Y=7056000
X3843 24 3805 ICV_1 $T=4608000 9840000 1 180 $X=4424000 $Y=9840000
X3844 24 3806 ICV_1 $T=4640000 5432000 1 180 $X=4456000 $Y=5432000
X3845 24 3807 ICV_1 $T=4656000 11232000 1 180 $X=4472000 $Y=11232000
X3846 24 3808 ICV_1 $T=4704000 4504000 1 180 $X=4520000 $Y=4504000
X3847 24 3809 ICV_1 $T=4736000 4736000 1 180 $X=4552000 $Y=4736000
X3848 24 3810 ICV_1 $T=4776000 7984000 1 180 $X=4592000 $Y=7984000
X3849 24 3811 ICV_1 $T=4920000 1952000 1 180 $X=4736000 $Y=1952000
X3850 24 3812 ICV_1 $T=4920000 7752000 1 180 $X=4736000 $Y=7752000
X3851 24 3813 ICV_1 $T=4936000 11000000 1 180 $X=4752000 $Y=11000000
X3852 24 3814 ICV_1 $T=4952000 4504000 1 180 $X=4768000 $Y=4504000
X3853 24 3815 ICV_1 $T=5104000 10072000 1 180 $X=4920000 $Y=10072000
X3854 24 3816 ICV_1 $T=5112000 1256000 1 180 $X=4928000 $Y=1256000
X3855 24 3817 ICV_1 $T=5128000 4736000 1 180 $X=4944000 $Y=4736000
X3856 24 3818 ICV_1 $T=5136000 4968000 1 180 $X=4952000 $Y=4968000
X3857 24 3819 ICV_1 $T=5176000 9144000 1 180 $X=4992000 $Y=9144000
X3858 24 3820 ICV_1 $T=5192000 5664000 1 180 $X=5008000 $Y=5664000
X3859 24 3821 ICV_1 $T=5192000 5896000 1 180 $X=5008000 $Y=5896000
X3860 24 3822 ICV_1 $T=5216000 9840000 1 180 $X=5032000 $Y=9840000
X3861 24 3823 ICV_1 $T=5280000 13088000 1 180 $X=5096000 $Y=13088000
X3862 24 3824 ICV_1 $T=5296000 5432000 1 180 $X=5112000 $Y=5432000
X3863 24 3825 ICV_1 $T=5304000 6128000 1 180 $X=5120000 $Y=6128000
X3864 24 3826 ICV_1 $T=5312000 8680000 1 180 $X=5128000 $Y=8680000
X3865 24 3827 ICV_1 $T=5328000 13320000 1 180 $X=5144000 $Y=13320000
X3866 24 3828 ICV_1 $T=5336000 1024000 1 180 $X=5152000 $Y=1024000
X3867 24 3829 ICV_1 $T=5352000 8216000 1 180 $X=5168000 $Y=8216000
X3868 24 3830 ICV_1 $T=5392000 6360000 1 180 $X=5208000 $Y=6360000
X3869 24 3831 ICV_1 $T=5424000 1256000 1 180 $X=5240000 $Y=1256000
X3870 24 3832 ICV_1 $T=5456000 9144000 1 180 $X=5272000 $Y=9144000
X3871 24 3833 ICV_1 $T=5504000 5200000 1 180 $X=5320000 $Y=5200000
X3872 24 3834 ICV_1 $T=5512000 12856000 1 180 $X=5328000 $Y=12856000
X3873 24 3835 ICV_1 $T=5536000 9376000 1 180 $X=5352000 $Y=9376000
X3874 24 3836 ICV_1 $T=5544000 5432000 1 180 $X=5360000 $Y=5432000
X3875 24 3837 ICV_1 $T=5552000 6128000 1 180 $X=5368000 $Y=6128000
X3876 24 3838 ICV_1 $T=5552000 7984000 1 180 $X=5368000 $Y=7984000
X3877 24 3839 ICV_1 $T=5672000 9608000 1 180 $X=5488000 $Y=9608000
X3878 24 3840 ICV_1 $T=5688000 4968000 1 180 $X=5504000 $Y=4968000
X3879 24 3841 ICV_1 $T=5696000 4504000 1 180 $X=5512000 $Y=4504000
X3880 24 3842 ICV_1 $T=5696000 6360000 1 180 $X=5512000 $Y=6360000
X3881 24 3843 ICV_1 $T=5704000 9144000 1 180 $X=5520000 $Y=9144000
X3882 24 3844 ICV_1 $T=5752000 6824000 1 180 $X=5568000 $Y=6824000
X3883 24 3845 ICV_1 $T=5776000 5664000 1 180 $X=5592000 $Y=5664000
X3884 24 3846 ICV_1 $T=5808000 5896000 1 180 $X=5624000 $Y=5896000
X3885 24 3847 ICV_1 $T=5816000 4736000 1 180 $X=5632000 $Y=4736000
X3886 24 3848 ICV_1 $T=5840000 7520000 1 180 $X=5656000 $Y=7520000
X3887 24 3849 ICV_1 $T=5880000 7056000 1 180 $X=5696000 $Y=7056000
X3888 24 3850 ICV_1 $T=5904000 792000 1 180 $X=5720000 $Y=792000
X3889 24 3851 ICV_1 $T=5936000 4968000 1 180 $X=5752000 $Y=4968000
X3890 24 3852 ICV_1 $T=5968000 9608000 1 180 $X=5784000 $Y=9608000
X3891 24 3853 ICV_1 $T=6056000 5896000 1 180 $X=5872000 $Y=5896000
X3892 24 3854 ICV_1 $T=6072000 6592000 1 180 $X=5888000 $Y=6592000
X3893 24 3855 ICV_1 $T=6080000 5664000 1 180 $X=5896000 $Y=5664000
X3894 24 3856 ICV_1 $T=6080000 6128000 1 180 $X=5896000 $Y=6128000
X3895 24 3857 ICV_1 $T=6184000 4968000 1 180 $X=6000000 $Y=4968000
X3896 24 3858 ICV_1 $T=6200000 4040000 1 180 $X=6016000 $Y=4040000
X3897 24 3859 ICV_1 $T=6216000 5200000 1 180 $X=6032000 $Y=5200000
X3898 24 3860 ICV_1 $T=6232000 4272000 1 180 $X=6048000 $Y=4272000
X3899 24 3861 ICV_1 $T=6256000 13320000 1 180 $X=6072000 $Y=13320000
X3900 24 3862 ICV_1 $T=6264000 12856000 1 180 $X=6080000 $Y=12856000
X3901 24 3863 ICV_1 $T=6304000 5896000 1 180 $X=6120000 $Y=5896000
X3902 24 3864 ICV_1 $T=6320000 6592000 1 180 $X=6136000 $Y=6592000
X3903 24 3865 ICV_1 $T=6328000 5664000 1 180 $X=6144000 $Y=5664000
X3904 24 3866 ICV_1 $T=6328000 6128000 1 180 $X=6144000 $Y=6128000
X3905 24 3867 ICV_1 $T=6328000 9608000 1 180 $X=6144000 $Y=9608000
X3906 24 3868 ICV_1 $T=6336000 6824000 1 180 $X=6152000 $Y=6824000
X3907 24 3869 ICV_1 $T=6360000 7752000 1 180 $X=6176000 $Y=7752000
X3908 24 3870 ICV_1 $T=6376000 9376000 1 180 $X=6192000 $Y=9376000
X3909 24 3871 ICV_1 $T=6400000 3112000 1 180 $X=6216000 $Y=3112000
X3910 24 3872 ICV_1 $T=6464000 5200000 1 180 $X=6280000 $Y=5200000
X3911 24 3873 ICV_1 $T=6480000 2648000 1 180 $X=6296000 $Y=2648000
X3912 24 3874 ICV_1 $T=6552000 5896000 1 180 $X=6368000 $Y=5896000
X3913 24 3875 ICV_1 $T=6560000 96000 1 180 $X=6376000 $Y=96000
X3914 24 3876 ICV_1 $T=6568000 6360000 1 180 $X=6384000 $Y=6360000
X3915 24 3877 ICV_1 $T=6576000 5664000 1 180 $X=6392000 $Y=5664000
X3916 24 3878 ICV_1 $T=6784000 7056000 1 180 $X=6600000 $Y=7056000
X3917 24 3879 ICV_1 $T=6808000 2184000 1 180 $X=6624000 $Y=2184000
X3918 24 3880 ICV_1 $T=6832000 6824000 1 180 $X=6648000 $Y=6824000
X3919 24 3881 ICV_1 $T=6872000 6592000 1 180 $X=6688000 $Y=6592000
X3920 24 3882 ICV_1 $T=6896000 5896000 1 180 $X=6712000 $Y=5896000
X3921 24 3883 ICV_1 $T=6912000 6360000 1 180 $X=6728000 $Y=6360000
X3922 24 3884 ICV_1 $T=6952000 3112000 1 180 $X=6768000 $Y=3112000
X3923 24 3885 ICV_1 $T=6960000 2648000 1 180 $X=6776000 $Y=2648000
X3924 24 3886 ICV_1 $T=6960000 11928000 1 180 $X=6776000 $Y=11928000
X3925 24 3887 ICV_1 $T=6992000 9376000 1 180 $X=6808000 $Y=9376000
X3926 24 3888 ICV_1 $T=7104000 1488000 1 180 $X=6920000 $Y=1488000
X3927 24 3889 ICV_1 $T=7120000 6592000 1 180 $X=6936000 $Y=6592000
X3928 24 3890 ICV_1 $T=7128000 9608000 1 180 $X=6944000 $Y=9608000
X3929 24 3891 ICV_1 $T=7144000 96000 1 180 $X=6960000 $Y=96000
X3930 24 3892 ICV_1 $T=7176000 11232000 1 180 $X=6992000 $Y=11232000
X3931 24 3893 ICV_1 $T=7200000 4968000 1 180 $X=7016000 $Y=4968000
X3932 24 3894 ICV_1 $T=7208000 792000 1 180 $X=7024000 $Y=792000
X3933 24 3895 ICV_1 $T=7208000 1256000 1 180 $X=7024000 $Y=1256000
X3934 24 3896 ICV_1 $T=7216000 560000 1 180 $X=7032000 $Y=560000
X3935 24 3897 ICV_1 $T=7224000 4272000 1 180 $X=7040000 $Y=4272000
X3936 24 3898 ICV_1 $T=7240000 9144000 1 180 $X=7056000 $Y=9144000
X3937 24 3899 ICV_1 $T=7240000 11464000 1 180 $X=7056000 $Y=11464000
X3938 24 3900 ICV_1 $T=7240000 11696000 1 180 $X=7056000 $Y=11696000
X3939 24 3901 ICV_1 $T=7240000 11928000 1 180 $X=7056000 $Y=11928000
X3940 24 3902 ICV_1 $T=7288000 9840000 1 180 $X=7104000 $Y=9840000
X3941 24 3903 ICV_1 $T=7344000 7288000 1 180 $X=7160000 $Y=7288000
X3942 24 3904 ICV_1 $T=7368000 328000 1 180 $X=7184000 $Y=328000
X3943 24 3905 ICV_1 $T=7424000 96000 1 180 $X=7240000 $Y=96000
X3944 24 3906 ICV_1 $T=7440000 9376000 1 180 $X=7256000 $Y=9376000
X3945 24 3907 ICV_1 $T=7448000 12160000 1 180 $X=7264000 $Y=12160000
X3946 24 3908 ICV_1 $T=7456000 792000 1 180 $X=7272000 $Y=792000
X3947 24 3909 ICV_1 $T=7472000 4272000 1 180 $X=7288000 $Y=4272000
X3948 24 3910 ICV_1 $T=7496000 2880000 1 180 $X=7312000 $Y=2880000
X3949 24 3911 ICV_1 $T=7504000 1720000 1 180 $X=7320000 $Y=1720000
X3950 24 3912 ICV_1 $T=7504000 10072000 1 180 $X=7320000 $Y=10072000
X3951 24 3913 ICV_1 $T=7528000 4736000 1 180 $X=7344000 $Y=4736000
X3952 24 3914 ICV_1 $T=7528000 9144000 1 180 $X=7344000 $Y=9144000
X3953 24 3915 ICV_1 $T=7528000 13320000 1 180 $X=7344000 $Y=13320000
X3954 24 3916 ICV_1 $T=7552000 8680000 1 180 $X=7368000 $Y=8680000
X3955 24 3917 ICV_1 $T=7568000 1952000 1 180 $X=7384000 $Y=1952000
X3956 24 3918 ICV_1 $T=7568000 3808000 1 180 $X=7384000 $Y=3808000
X3957 24 3919 ICV_1 $T=7592000 7520000 1 180 $X=7408000 $Y=7520000
X3958 24 3920 ICV_1 $T=7608000 6824000 1 180 $X=7424000 $Y=6824000
X3959 24 3921 ICV_1 $T=7608000 7056000 1 180 $X=7424000 $Y=7056000
X3960 24 3922 ICV_1 $T=7640000 6128000 1 180 $X=7456000 $Y=6128000
X3961 24 3923 ICV_1 $T=7640000 12624000 1 180 $X=7456000 $Y=12624000
X3962 24 3924 ICV_1 $T=7648000 12392000 1 180 $X=7464000 $Y=12392000
X3963 24 3925 ICV_1 $T=7664000 2184000 1 180 $X=7480000 $Y=2184000
X3964 24 3926 ICV_1 $T=7680000 4040000 1 180 $X=7496000 $Y=4040000
X3965 24 3927 ICV_1 $T=7688000 11928000 1 180 $X=7504000 $Y=11928000
X3966 24 3928 ICV_1 $T=7776000 13552000 1 180 $X=7592000 $Y=13552000
X3967 24 3929 ICV_1 $T=7816000 1256000 1 180 $X=7632000 $Y=1256000
X3968 24 3930 ICV_1 $T=7816000 2648000 1 180 $X=7632000 $Y=2648000
X3969 24 3931 ICV_1 $T=7824000 1024000 1 180 $X=7640000 $Y=1024000
X3970 24 3932 ICV_1 $T=7856000 2880000 1 180 $X=7672000 $Y=2880000
X3971 24 3933 ICV_1 $T=7872000 1488000 1 180 $X=7688000 $Y=1488000
X3972 24 3934 ICV_1 $T=7888000 12624000 1 180 $X=7704000 $Y=12624000
X3973 24 3935 ICV_1 $T=7896000 7520000 1 180 $X=7712000 $Y=7520000
X3974 24 3936 ICV_1 $T=8072000 1024000 1 180 $X=7888000 $Y=1024000
X3975 24 3937 ICV_1 $T=8160000 2184000 1 180 $X=7976000 $Y=2184000
X3976 24 3938 ICV_1 $T=8216000 2416000 1 180 $X=8032000 $Y=2416000
X3977 24 3939 ICV_1 $T=8256000 12856000 1 180 $X=8072000 $Y=12856000
X3978 24 3940 ICV_1 $T=8264000 7288000 1 180 $X=8080000 $Y=7288000
X3979 24 3941 ICV_1 $T=8272000 5896000 1 180 $X=8088000 $Y=5896000
X3980 24 3942 ICV_1 $T=8304000 7752000 1 180 $X=8120000 $Y=7752000
X3981 24 3943 ICV_1 $T=8368000 2648000 1 180 $X=8184000 $Y=2648000
X3982 24 3944 ICV_1 $T=8368000 4040000 1 180 $X=8184000 $Y=4040000
X3983 24 3945 ICV_1 $T=8368000 10304000 1 180 $X=8184000 $Y=10304000
X3984 24 3946 ICV_1 $T=8408000 2184000 1 180 $X=8224000 $Y=2184000
X3985 24 3947 ICV_1 $T=8424000 12160000 1 180 $X=8240000 $Y=12160000
X3986 24 3948 ICV_1 $T=8504000 12856000 1 180 $X=8320000 $Y=12856000
X3987 24 3949 ICV_1 $T=8512000 7288000 1 180 $X=8328000 $Y=7288000
X3988 24 3950 ICV_1 $T=8512000 9840000 1 180 $X=8328000 $Y=9840000
X3989 24 3951 ICV_1 $T=8520000 5896000 1 180 $X=8336000 $Y=5896000
X3990 24 3952 ICV_1 $T=8536000 11000000 1 180 $X=8352000 $Y=11000000
X3991 24 3953 ICV_1 $T=8552000 7984000 1 180 $X=8368000 $Y=7984000
X3992 24 3954 ICV_1 $T=8560000 10072000 1 180 $X=8376000 $Y=10072000
X3993 24 3955 ICV_1 $T=8560000 13552000 1 180 $X=8376000 $Y=13552000
X3994 24 3956 ICV_1 $T=8576000 12624000 1 180 $X=8392000 $Y=12624000
X3995 24 3957 ICV_1 $T=8600000 13320000 1 180 $X=8416000 $Y=13320000
X3996 24 3958 ICV_1 $T=8616000 4040000 1 180 $X=8432000 $Y=4040000
X3997 24 3959 ICV_1 $T=8640000 2416000 1 180 $X=8456000 $Y=2416000
X3998 24 3960 ICV_1 $T=8648000 12392000 1 180 $X=8464000 $Y=12392000
X3999 24 3961 ICV_1 $T=8656000 2184000 1 180 $X=8472000 $Y=2184000
X4000 24 3962 ICV_1 $T=8664000 1952000 1 180 $X=8480000 $Y=1952000
X4001 24 3963 ICV_1 $T=8664000 3808000 1 180 $X=8480000 $Y=3808000
X4002 24 3964 ICV_1 $T=8680000 3112000 1 180 $X=8496000 $Y=3112000
X4003 24 3965 ICV_1 $T=8696000 9376000 1 180 $X=8512000 $Y=9376000
X4004 24 3966 ICV_1 $T=8704000 2880000 1 180 $X=8520000 $Y=2880000
X4005 24 3967 ICV_1 $T=8704000 12160000 1 180 $X=8520000 $Y=12160000
X4006 24 3968 ICV_1 $T=8712000 9608000 1 180 $X=8528000 $Y=9608000
X4007 24 3969 ICV_1 $T=8760000 13088000 1 180 $X=8576000 $Y=13088000
X4008 24 3970 ICV_1 $T=8808000 13552000 1 180 $X=8624000 $Y=13552000
X4009 24 3971 ICV_1 $T=8824000 12624000 1 180 $X=8640000 $Y=12624000
X4010 24 3972 ICV_1 $T=8832000 7984000 1 180 $X=8648000 $Y=7984000
X4011 24 3973 ICV_1 $T=8872000 1024000 1 180 $X=8688000 $Y=1024000
X4012 24 3974 ICV_1 $T=8888000 2416000 1 180 $X=8704000 $Y=2416000
X4013 24 3975 ICV_1 $T=8896000 12392000 1 180 $X=8712000 $Y=12392000
X4014 24 3976 ICV_1 $T=8904000 2184000 1 180 $X=8720000 $Y=2184000
X4015 24 3977 ICV_1 $T=8928000 3112000 1 180 $X=8744000 $Y=3112000
X4016 24 3978 ICV_1 $T=8952000 2880000 1 180 $X=8768000 $Y=2880000
X4017 24 3979 ICV_1 $T=8960000 9144000 1 180 $X=8776000 $Y=9144000
X4018 24 3980 ICV_1 $T=9008000 1952000 1 180 $X=8824000 $Y=1952000
X4019 24 3981 ICV_1 $T=9032000 3576000 1 180 $X=8848000 $Y=3576000
X4020 24 3982 ICV_1 $T=9048000 8216000 1 180 $X=8864000 $Y=8216000
X4021 24 3983 ICV_1 $T=9056000 8448000 1 180 $X=8872000 $Y=8448000
X4022 24 3984 ICV_1 $T=9056000 13552000 1 180 $X=8872000 $Y=13552000
X4023 24 3985 ICV_1 $T=9064000 13088000 1 180 $X=8880000 $Y=13088000
X4024 24 3986 ICV_1 $T=9136000 13320000 1 180 $X=8952000 $Y=13320000
X4025 24 3987 ICV_1 $T=9144000 2648000 1 180 $X=8960000 $Y=2648000
X4026 24 3988 ICV_1 $T=9256000 6824000 1 180 $X=9072000 $Y=6824000
X4027 24 3989 ICV_1 $T=9272000 8680000 1 180 $X=9088000 $Y=8680000
X4028 24 3990 ICV_1 $T=9280000 12624000 1 180 $X=9096000 $Y=12624000
X4029 24 3991 ICV_1 $T=9304000 13552000 1 180 $X=9120000 $Y=13552000
X4030 24 3992 ICV_1 $T=9312000 13088000 1 180 $X=9128000 $Y=13088000
X4031 24 3993 ICV_1 $T=9368000 12392000 1 180 $X=9184000 $Y=12392000
X4032 24 3994 ICV_1 $T=9392000 2648000 1 180 $X=9208000 $Y=2648000
X4033 24 3995 ICV_1 $T=9416000 792000 1 180 $X=9232000 $Y=792000
X4034 24 3996 ICV_1 $T=9416000 1024000 1 180 $X=9232000 $Y=1024000
X4035 24 3997 ICV_1 $T=9424000 12160000 1 180 $X=9240000 $Y=12160000
X4036 24 3998 ICV_1 $T=9440000 96000 1 180 $X=9256000 $Y=96000
X4037 24 3999 ICV_1 $T=9440000 3808000 1 180 $X=9256000 $Y=3808000
X4038 24 4000 ICV_1 $T=9448000 13320000 1 180 $X=9264000 $Y=13320000
X4039 24 4001 ICV_1 $T=9520000 7520000 1 180 $X=9336000 $Y=7520000
X4040 24 4002 ICV_1 $T=9520000 8680000 1 180 $X=9336000 $Y=8680000
X4041 24 4003 ICV_1 $T=9536000 560000 1 180 $X=9352000 $Y=560000
X4042 24 4004 ICV_1 $T=9600000 7984000 1 180 $X=9416000 $Y=7984000
X4043 24 4005 ICV_1 $T=9608000 7288000 1 180 $X=9424000 $Y=7288000
X4044 24 4006 ICV_1 $T=9632000 13552000 1 180 $X=9448000 $Y=13552000
X4045 24 4007 ICV_1 $T=9664000 1024000 1 180 $X=9480000 $Y=1024000
X4046 24 4008 ICV_1 $T=9672000 9608000 1 180 $X=9488000 $Y=9608000
X4047 24 4009 ICV_1 $T=9696000 13320000 1 180 $X=9512000 $Y=13320000
X4048 24 4010 ICV_1 $T=9728000 4968000 1 180 $X=9544000 $Y=4968000
X4049 24 4011 ICV_1 $T=9736000 9376000 1 180 $X=9552000 $Y=9376000
X4050 24 4012 ICV_1 $T=9776000 792000 1 180 $X=9592000 $Y=792000
X4051 24 4013 ICV_1 $T=9776000 4272000 1 180 $X=9592000 $Y=4272000
X4052 24 4014 ICV_1 $T=9776000 8912000 1 180 $X=9592000 $Y=8912000
X4053 24 4015 ICV_1 $T=9808000 12160000 1 180 $X=9624000 $Y=12160000
X4054 24 4016 ICV_1 $T=9832000 4504000 1 180 $X=9648000 $Y=4504000
X4055 24 4017 ICV_1 $T=9872000 5432000 1 180 $X=9688000 $Y=5432000
X4056 24 4018 ICV_1 $T=9928000 4040000 1 180 $X=9744000 $Y=4040000
X4057 24 4019 ICV_1 $T=9976000 4968000 1 180 $X=9792000 $Y=4968000
X4058 24 4020 ICV_1 $T=9984000 9376000 1 180 $X=9800000 $Y=9376000
X4059 24 4021 ICV_1 $T=10024000 792000 1 180 $X=9840000 $Y=792000
X4060 24 4022 ICV_1 $T=10048000 8448000 1 180 $X=9864000 $Y=8448000
X4061 24 4023 ICV_1 $T=10056000 5200000 1 180 $X=9872000 $Y=5200000
X4062 24 4024 ICV_1 $T=10064000 2184000 1 180 $X=9880000 $Y=2184000
X4063 24 4025 ICV_1 $T=10104000 8912000 1 180 $X=9920000 $Y=8912000
X4064 24 4026 ICV_1 $T=10176000 11000000 1 180 $X=9992000 $Y=11000000
X4065 24 4027 ICV_1 $T=10184000 1256000 1 180 $X=10000000 $Y=1256000
X4066 24 4028 ICV_1 $T=10240000 10536000 1 180 $X=10056000 $Y=10536000
X4067 24 4029 ICV_1 $T=10272000 792000 1 180 $X=10088000 $Y=792000
X4068 24 4030 ICV_1 $T=10280000 9608000 1 180 $X=10096000 $Y=9608000
X4069 24 4031 ICV_1 $T=10288000 4040000 1 180 $X=10104000 $Y=4040000
X4070 24 4032 ICV_1 $T=10296000 5896000 1 180 $X=10112000 $Y=5896000
X4071 24 4033 ICV_1 $T=10312000 2184000 1 180 $X=10128000 $Y=2184000
X4072 24 4034 ICV_1 $T=10328000 1024000 1 180 $X=10144000 $Y=1024000
X4073 24 4035 ICV_1 $T=10336000 560000 1 180 $X=10152000 $Y=560000
X4074 24 4036 ICV_1 $T=10392000 5200000 1 180 $X=10208000 $Y=5200000
X4075 24 4037 ICV_1 $T=10464000 1256000 1 180 $X=10280000 $Y=1256000
X4076 24 4038 ICV_1 $T=10504000 7984000 1 180 $X=10320000 $Y=7984000
X4077 24 4039 ICV_1 $T=10536000 4040000 1 180 $X=10352000 $Y=4040000
X4078 24 4040 ICV_1 $T=10552000 4272000 1 180 $X=10368000 $Y=4272000
X4079 24 4041 ICV_1 $T=10616000 6592000 1 180 $X=10432000 $Y=6592000
X4080 24 4042 ICV_1 $T=10616000 9144000 1 180 $X=10432000 $Y=9144000
X4081 24 4043 ICV_1 $T=10656000 1952000 1 180 $X=10472000 $Y=1952000
X4082 24 4044 ICV_1 $T=10664000 2648000 1 180 $X=10480000 $Y=2648000
X4083 24 4045 ICV_1 $T=10704000 11232000 1 180 $X=10520000 $Y=11232000
X4084 24 4046 ICV_1 $T=10728000 1720000 1 180 $X=10544000 $Y=1720000
X4085 24 4047 ICV_1 $T=10736000 2880000 1 180 $X=10552000 $Y=2880000
X4086 24 4048 ICV_1 $T=10744000 9376000 1 180 $X=10560000 $Y=9376000
X4087 24 4049 ICV_1 $T=10784000 7056000 1 180 $X=10600000 $Y=7056000
X4088 24 4050 ICV_1 $T=10824000 11464000 1 180 $X=10640000 $Y=11464000
X4089 24 4051 ICV_1 $T=10864000 9144000 1 180 $X=10680000 $Y=9144000
X4090 24 4052 ICV_1 $T=10880000 8912000 1 180 $X=10696000 $Y=8912000
X4091 24 4053 ICV_1 $T=10912000 2648000 1 180 $X=10728000 $Y=2648000
X4092 24 4054 ICV_1 $T=10936000 1952000 1 180 $X=10752000 $Y=1952000
X4093 24 4055 ICV_1 $T=10976000 1720000 1 180 $X=10792000 $Y=1720000
X4094 24 4056 ICV_1 $T=10984000 2880000 1 180 $X=10800000 $Y=2880000
X4095 24 4057 ICV_1 $T=11112000 11464000 1 180 $X=10928000 $Y=11464000
X4096 24 4058 ICV_1 $T=11176000 9144000 1 180 $X=10992000 $Y=9144000
X4097 24 4059 ICV_1 $T=11344000 10304000 1 180 $X=11160000 $Y=10304000
X4098 24 4060 ICV_1 $T=11392000 10072000 1 180 $X=11208000 $Y=10072000
X4099 24 4061 ICV_1 $T=11424000 11464000 1 180 $X=11240000 $Y=11464000
X4100 24 4062 ICV_1 $T=11432000 11000000 1 180 $X=11248000 $Y=11000000
X4101 24 4063 ICV_1 $T=11464000 5664000 1 180 $X=11280000 $Y=5664000
X4102 24 4064 ICV_1 $T=11480000 13088000 1 180 $X=11296000 $Y=13088000
X4103 24 4065 ICV_1 $T=11488000 12856000 1 180 $X=11304000 $Y=12856000
X4104 24 4066 ICV_1 $T=11536000 9144000 1 180 $X=11352000 $Y=9144000
X4105 24 4067 ICV_1 $T=11536000 9376000 1 180 $X=11352000 $Y=9376000
X4106 24 4068 ICV_1 $T=11536000 10768000 1 180 $X=11352000 $Y=10768000
X4107 24 4069 ICV_1 $T=11584000 5896000 1 180 $X=11400000 $Y=5896000
X4108 24 4070 ICV_1 $T=11712000 5664000 1 180 $X=11528000 $Y=5664000
X4109 24 4071 ICV_1 $T=11736000 3344000 1 180 $X=11552000 $Y=3344000
X4110 24 4072 ICV_1 $T=11736000 3576000 1 180 $X=11552000 $Y=3576000
X4111 24 4073 ICV_1 $T=11752000 5432000 1 180 $X=11568000 $Y=5432000
X4112 24 4074 ICV_1 $T=11832000 10072000 1 180 $X=11648000 $Y=10072000
X4113 24 4075 ICV_1 $T=11912000 2184000 1 180 $X=11728000 $Y=2184000
X4114 24 4076 ICV_1 $T=11952000 7984000 1 180 $X=11768000 $Y=7984000
X4115 24 4077 ICV_1 $T=11960000 5664000 1 180 $X=11776000 $Y=5664000
X4116 24 4078 ICV_1 $T=11968000 10304000 1 180 $X=11784000 $Y=10304000
X4117 24 4079 ICV_1 $T=12032000 5432000 1 180 $X=11848000 $Y=5432000
X4118 24 4080 ICV_1 $T=12032000 8216000 1 180 $X=11848000 $Y=8216000
X4119 24 4081 ICV_1 $T=12032000 9144000 1 180 $X=11848000 $Y=9144000
X4120 24 4082 ICV_1 $T=12032000 10536000 1 180 $X=11848000 $Y=10536000
X4121 24 4083 ICV_1 $T=12160000 10072000 1 180 $X=11976000 $Y=10072000
X4122 24 4084 ICV_1 $T=12200000 7984000 1 180 $X=12016000 $Y=7984000
X4123 24 4085 ICV_1 $T=12200000 11232000 1 180 $X=12016000 $Y=11232000
X4124 24 4086 ICV_1 $T=12208000 5664000 1 180 $X=12024000 $Y=5664000
X4125 24 4087 ICV_1 $T=12208000 5896000 1 180 $X=12024000 $Y=5896000
X4126 24 4088 ICV_1 $T=12216000 6128000 1 180 $X=12032000 $Y=6128000
X4127 24 4089 ICV_1 $T=12216000 6592000 1 180 $X=12032000 $Y=6592000
X4128 24 4090 ICV_1 $T=12216000 9376000 1 180 $X=12032000 $Y=9376000
X4129 24 4091 ICV_1 $T=12216000 9608000 1 180 $X=12032000 $Y=9608000
X4130 24 4092 ICV_1 $T=12216000 9840000 1 180 $X=12032000 $Y=9840000
X4131 24 4093 ICV_1 $T=12216000 10304000 1 180 $X=12032000 $Y=10304000
X4132 24 4094 ICV_1 $T=12280000 6360000 1 180 $X=12096000 $Y=6360000
X4133 24 4095 ICV_1 $T=12280000 9144000 1 180 $X=12096000 $Y=9144000
X4134 24 4096 ICV_1 $T=12360000 8680000 1 180 $X=12176000 $Y=8680000
X4135 24 4082 ICV_2 $T=11664000 10536000 1 180 $X=11480000 $Y=10536000
X4136 24 4097 ICV_2 $T=11952000 13320000 1 180 $X=11768000 $Y=13320000
X4137 24 4097 ICV_2 $T=12320000 13320000 1 180 $X=12136000 $Y=13320000
X4138 24 4098 ICV_2 $T=12344000 13552000 1 180 $X=12160000 $Y=13552000
X4139 24 ICV_3 $T=10176000 96000 0 0 $X=10176000 $Y=96000
X4140 24 ICV_3 $T=11680000 8680000 0 0 $X=11680000 $Y=8680000
X4141 24 ICV_3 $T=11872000 1720000 0 0 $X=11872000 $Y=1720000
X4142 24 ICV_3 $T=12160000 6824000 0 0 $X=12160000 $Y=6824000
X4143 24 2508 ICV_4 $T=624000 12624000 0 0 $X=624000 $Y=12624000
X4144 24 2681 ICV_4 $T=4056000 10536000 0 0 $X=4056000 $Y=10536000
X4145 24 443 ICV_4 $T=4104000 5896000 0 0 $X=4104000 $Y=5896000
X4146 24 485 ICV_4 $T=4536000 11928000 0 0 $X=4536000 $Y=11928000
X4147 24 3819 ICV_4 $T=4624000 9144000 0 0 $X=4624000 $Y=9144000
X4148 24 4099 ICV_4 $T=6536000 10304000 0 0 $X=6536000 $Y=10304000
X4149 24 2344 ICV_4 $T=8184000 4736000 0 0 $X=8184000 $Y=4736000
X4150 24 4100 ICV_4 $T=8552000 11464000 0 0 $X=8552000 $Y=11464000
X4151 24 824 ICV_4 $T=8632000 11232000 0 0 $X=8632000 $Y=11232000
X4152 24 3995 ICV_4 $T=8864000 792000 0 0 $X=8864000 $Y=792000
X4153 24 851 ICV_4 $T=9224000 3576000 0 0 $X=9224000 $Y=3576000
X4154 24 2352 ICV_4 $T=9664000 5664000 0 0 $X=9664000 $Y=5664000
X4155 24 2866 ICV_4 $T=10016000 11464000 0 0 $X=10016000 $Y=11464000
X4156 24 4101 ICV_4 $T=10392000 7752000 0 0 $X=10392000 $Y=7752000
X4157 24 4102 ICV_4 $T=10672000 11928000 0 0 $X=10672000 $Y=11928000
X4158 24 4103 ICV_4 $T=10888000 3344000 0 0 $X=10888000 $Y=3344000
X4159 24 967 ICV_4 $T=11360000 2880000 0 0 $X=11360000 $Y=2880000
X4160 24 4104 ICV_4 $T=12160000 2880000 0 0 $X=12160000 $Y=2880000
X4161 24 4105 ICV_4 $T=12160000 3576000 0 0 $X=12160000 $Y=3576000
X4162 24 4106 ICV_4 $T=12160000 4504000 0 0 $X=12160000 $Y=4504000
X4163 24 4107 nand04 $T=648000 7520000 0 0 $X=648000 $Y=7520000
X4164 24 4108 nand04 $T=760000 6128000 0 0 $X=760000 $Y=6128000
X4165 24 4109 nand04 $T=849000 11928000 1 180 $X=800000 $Y=11928000
X4166 24 4110 nand04 $T=865000 11232000 1 180 $X=816000 $Y=11232000
X4167 24 4111 nand04 $T=905000 5432000 1 180 $X=856000 $Y=5432000
X4168 24 4112 nand04 $T=872000 13088000 0 0 $X=872000 $Y=13088000
X4169 24 4113 nand04 $T=961000 3808000 1 180 $X=912000 $Y=3808000
X4170 24 4114 nand04 $T=977000 11232000 1 180 $X=928000 $Y=11232000
X4171 24 4115 nand04 $T=928000 13088000 0 0 $X=928000 $Y=13088000
X4172 24 4116 nand04 $T=1001000 11928000 1 180 $X=952000 $Y=11928000
X4173 24 4117 nand04 $T=1112000 7288000 0 0 $X=1112000 $Y=7288000
X4174 24 4118 nand04 $T=1120000 4736000 0 0 $X=1120000 $Y=4736000
X4175 24 4119 nand04 $T=1128000 6128000 0 0 $X=1128000 $Y=6128000
X4176 24 4120 nand04 $T=1209000 12856000 1 180 $X=1160000 $Y=12856000
X4177 24 4121 nand04 $T=1233000 5432000 1 180 $X=1184000 $Y=5432000
X4178 24 4122 nand04 $T=1200000 7984000 0 0 $X=1200000 $Y=7984000
X4179 24 4123 nand04 $T=1200000 9144000 0 0 $X=1200000 $Y=9144000
X4180 24 4124 nand04 $T=1208000 4736000 0 0 $X=1208000 $Y=4736000
X4181 24 4125 nand04 $T=1256000 9144000 0 0 $X=1256000 $Y=9144000
X4182 24 4126 nand04 $T=1568000 7520000 0 0 $X=1568000 $Y=7520000
X4183 24 4127 nand04 $T=1632000 6128000 0 0 $X=1632000 $Y=6128000
X4184 24 4128 nand04 $T=1672000 2880000 0 0 $X=1672000 $Y=2880000
X4185 24 4129 nand04 $T=1801000 11232000 1 180 $X=1752000 $Y=11232000
X4186 24 4130 nand04 $T=1784000 9608000 0 0 $X=1784000 $Y=9608000
X4187 24 4131 nand04 $T=1841000 4736000 1 180 $X=1792000 $Y=4736000
X4188 24 4132 nand04 $T=1872000 7288000 0 0 $X=1872000 $Y=7288000
X4189 24 4133 nand04 $T=1880000 12392000 0 0 $X=1880000 $Y=12392000
X4190 24 4134 nand04 $T=1920000 7752000 0 0 $X=1920000 $Y=7752000
X4191 24 4135 nand04 $T=1976000 2416000 0 0 $X=1976000 $Y=2416000
X4192 24 4136 nand04 $T=2033000 13088000 1 180 $X=1984000 $Y=13088000
X4193 24 4137 nand04 $T=2048000 6128000 0 0 $X=2048000 $Y=6128000
X4194 24 4138 nand04 $T=2104000 4040000 0 0 $X=2104000 $Y=4040000
X4195 24 4139 nand04 $T=2192000 1952000 0 0 $X=2192000 $Y=1952000
X4196 24 4140 nand04 $T=2273000 9144000 1 180 $X=2224000 $Y=9144000
X4197 24 4141 nand04 $T=2272000 5896000 0 0 $X=2272000 $Y=5896000
X4198 24 4142 nand04 $T=2464000 11232000 0 0 $X=2464000 $Y=11232000
X4199 24 4143 nand04 $T=2472000 4504000 0 0 $X=2472000 $Y=4504000
X4200 24 4144 nand04 $T=2601000 9608000 1 180 $X=2552000 $Y=9608000
X4201 24 4145 nand04 $T=2576000 4504000 0 0 $X=2576000 $Y=4504000
X4202 24 4146 nand04 $T=2680000 7288000 0 0 $X=2680000 $Y=7288000
X4203 24 2308 nand04 $T=2704000 5664000 0 0 $X=2704000 $Y=5664000
X4204 24 4147 nand04 $T=2849000 12856000 1 180 $X=2800000 $Y=12856000
X4205 24 2309 nand04 $T=2865000 4504000 1 180 $X=2816000 $Y=4504000
X4206 24 4148 nand04 $T=2889000 9144000 1 180 $X=2840000 $Y=9144000
X4207 24 4149 nand04 $T=2961000 7984000 1 180 $X=2912000 $Y=7984000
X4208 24 4150 nand04 $T=3208000 11000000 0 0 $X=3208000 $Y=11000000
X4209 24 4151 nand04 $T=3320000 12856000 0 0 $X=3320000 $Y=12856000
X4210 24 4152 nand04 $T=3376000 9144000 0 0 $X=3376000 $Y=9144000
X4211 24 4153 nand04 $T=3513000 11464000 1 180 $X=3464000 $Y=11464000
X4212 24 4154 nand04 $T=3569000 9608000 1 180 $X=3520000 $Y=9608000
X4213 24 4155 nand04 $T=3560000 10768000 0 0 $X=3560000 $Y=10768000
X4214 24 4156 nand04 $T=3672000 5432000 0 0 $X=3672000 $Y=5432000
X4215 24 4157 nand04 $T=3721000 12160000 1 180 $X=3672000 $Y=12160000
X4216 24 4158 nand04 $T=3704000 4040000 0 0 $X=3704000 $Y=4040000
X4217 24 4159 nand04 $T=3785000 5664000 1 180 $X=3736000 $Y=5664000
X4218 24 4160 nand04 $T=3736000 6360000 0 0 $X=3736000 $Y=6360000
X4219 24 4161 nand04 $T=3809000 7752000 1 180 $X=3760000 $Y=7752000
X4220 24 4162 nand04 $T=3784000 4968000 0 0 $X=3784000 $Y=4968000
X4221 24 4163 nand04 $T=3792000 4504000 0 0 $X=3792000 $Y=4504000
X4222 24 4164 nand04 $T=3841000 12392000 1 180 $X=3792000 $Y=12392000
X4223 24 4165 nand04 $T=3865000 7752000 1 180 $X=3816000 $Y=7752000
X4224 24 4166 nand04 $T=3921000 5200000 1 180 $X=3872000 $Y=5200000
X4225 24 4167 nand04 $T=3936000 792000 0 0 $X=3936000 $Y=792000
X4226 24 4168 nand04 $T=4025000 9608000 1 180 $X=3976000 $Y=9608000
X4227 24 4169 nand04 $T=4000000 2184000 0 0 $X=4000000 $Y=2184000
X4228 24 4170 nand04 $T=4000000 12392000 0 0 $X=4000000 $Y=12392000
X4229 24 4171 nand04 $T=4024000 1952000 0 0 $X=4024000 $Y=1952000
X4230 24 4172 nand04 $T=4097000 7056000 1 180 $X=4048000 $Y=7056000
X4231 24 4173 nand04 $T=4097000 11696000 1 180 $X=4048000 $Y=11696000
X4232 24 4174 nand04 $T=4129000 7520000 1 180 $X=4080000 $Y=7520000
X4233 24 4175 nand04 $T=4249000 3344000 1 180 $X=4200000 $Y=3344000
X4234 24 4176 nand04 $T=4216000 8912000 0 0 $X=4216000 $Y=8912000
X4235 24 4177 nand04 $T=4224000 1024000 0 0 $X=4224000 $Y=1024000
X4236 24 4178 nand04 $T=4273000 11000000 1 180 $X=4224000 $Y=11000000
X4237 24 4179 nand04 $T=4320000 9144000 0 0 $X=4320000 $Y=9144000
X4238 24 4180 nand04 $T=4328000 9608000 0 0 $X=4328000 $Y=9608000
X4239 24 4181 nand04 $T=4441000 12856000 1 180 $X=4392000 $Y=12856000
X4240 24 4182 nand04 $T=4465000 11232000 1 180 $X=4416000 $Y=11232000
X4241 24 4183 nand04 $T=4545000 4736000 1 180 $X=4496000 $Y=4736000
X4242 24 4184 nand04 $T=4729000 7288000 1 180 $X=4680000 $Y=7288000
X4243 24 4185 nand04 $T=4745000 792000 1 180 $X=4696000 $Y=792000
X4244 24 4186 nand04 $T=4712000 2184000 0 0 $X=4712000 $Y=2184000
X4245 24 4187 nand04 $T=4761000 5664000 1 180 $X=4712000 $Y=5664000
X4246 24 4188 nand04 $T=4808000 12392000 0 0 $X=4808000 $Y=12392000
X4247 24 4189 nand04 $T=4929000 5432000 1 180 $X=4880000 $Y=5432000
X4248 24 4190 nand04 $T=4896000 5664000 0 0 $X=4896000 $Y=5664000
X4249 24 4191 nand04 $T=4952000 6128000 0 0 $X=4952000 $Y=6128000
X4250 24 4192 nand04 $T=5025000 9840000 1 180 $X=4976000 $Y=9840000
X4251 24 4193 nand04 $T=4984000 7752000 0 0 $X=4984000 $Y=7752000
X4252 24 4194 nand04 $T=5049000 11000000 1 180 $X=5000000 $Y=11000000
X4253 24 4195 nand04 $T=5048000 2416000 0 0 $X=5048000 $Y=2416000
X4254 24 4196 nand04 $T=5064000 560000 0 0 $X=5064000 $Y=560000
X4255 24 4197 nand04 $T=5145000 6360000 1 180 $X=5096000 $Y=6360000
X4256 24 4198 nand04 $T=5104000 792000 0 0 $X=5104000 $Y=792000
X4257 24 4199 nand04 $T=5201000 8912000 1 180 $X=5152000 $Y=8912000
X4258 24 4200 nand04 $T=5176000 560000 0 0 $X=5176000 $Y=560000
X4259 24 4201 nand04 $T=5233000 11928000 1 180 $X=5184000 $Y=11928000
X4260 24 4202 nand04 $T=5265000 12856000 1 180 $X=5216000 $Y=12856000
X4261 24 4203 nand04 $T=5336000 4040000 0 0 $X=5336000 $Y=4040000
X4262 24 4204 nand04 $T=5481000 7752000 1 180 $X=5432000 $Y=7752000
X4263 24 4205 nand04 $T=5480000 5664000 0 0 $X=5480000 $Y=5664000
X4264 24 4206 nand04 $T=5488000 3576000 0 0 $X=5488000 $Y=3576000
X4265 24 4207 nand04 $T=5536000 6592000 0 0 $X=5536000 $Y=6592000
X4266 24 4208 nand04 $T=5585000 7288000 1 180 $X=5536000 $Y=7288000
X4267 24 4209 nand04 $T=5640000 10768000 0 0 $X=5640000 $Y=10768000
X4268 24 4210 nand04 $T=5881000 7288000 1 180 $X=5832000 $Y=7288000
X4269 24 4211 nand04 $T=5888000 2880000 0 0 $X=5888000 $Y=2880000
X4270 24 4212 nand04 $T=5928000 11696000 0 0 $X=5928000 $Y=11696000
X4271 24 4213 nand04 $T=5936000 2416000 0 0 $X=5936000 $Y=2416000
X4272 24 4214 nand04 $T=5968000 792000 0 0 $X=5968000 $Y=792000
X4273 24 4215 nand04 $T=5984000 12624000 0 0 $X=5984000 $Y=12624000
X4274 24 4216 nand04 $T=6032000 9376000 0 0 $X=6032000 $Y=9376000
X4275 24 4217 nand04 $T=6081000 9608000 1 180 $X=6032000 $Y=9608000
X4276 24 4218 nand04 $T=6145000 3808000 1 180 $X=6096000 $Y=3808000
X4277 24 4219 nand04 $T=6369000 9144000 1 180 $X=6320000 $Y=9144000
X4278 24 4220 nand04 $T=6584000 4736000 0 0 $X=6584000 $Y=4736000
X4279 24 4221 nand04 $T=6632000 3576000 0 0 $X=6632000 $Y=3576000
X4280 24 4222 nand04 $T=6713000 6128000 1 180 $X=6664000 $Y=6128000
X4281 24 4223 nand04 $T=6761000 2880000 1 180 $X=6712000 $Y=2880000
X4282 24 4224 nand04 $T=6744000 2416000 0 0 $X=6744000 $Y=2416000
X4283 24 4225 nand04 $T=6793000 13088000 1 180 $X=6744000 $Y=13088000
X4284 24 4226 nand04 $T=6792000 1024000 0 0 $X=6792000 $Y=1024000
X4285 24 4227 nand04 $T=6881000 6128000 1 180 $X=6832000 $Y=6128000
X4286 24 4228 nand04 $T=6832000 8912000 0 0 $X=6832000 $Y=8912000
X4287 24 4229 nand04 $T=6937000 328000 1 180 $X=6888000 $Y=328000
X4288 24 4230 nand04 $T=6928000 1024000 0 0 $X=6928000 $Y=1024000
X4289 24 4231 nand04 $T=6936000 11232000 0 0 $X=6936000 $Y=11232000
X4290 24 4232 nand04 $T=6992000 9840000 0 0 $X=6992000 $Y=9840000
X4291 24 4233 nand04 $T=7049000 4504000 1 180 $X=7000000 $Y=4504000
X4292 24 4234 nand04 $T=7000000 11696000 0 0 $X=7000000 $Y=11696000
X4293 24 4235 nand04 $T=7072000 7520000 0 0 $X=7072000 $Y=7520000
X4294 24 4236 nand04 $T=7129000 9376000 1 180 $X=7080000 $Y=9376000
X4295 24 4237 nand04 $T=7129000 12160000 1 180 $X=7080000 $Y=12160000
X4296 24 4238 nand04 $T=7273000 4504000 1 180 $X=7224000 $Y=4504000
X4297 24 4239 nand04 $T=7296000 7520000 0 0 $X=7296000 $Y=7520000
X4298 24 4240 nand04 $T=7336000 1024000 0 0 $X=7336000 $Y=1024000
X4299 24 4241 nand04 $T=7401000 12392000 1 180 $X=7352000 $Y=12392000
X4300 24 4242 nand04 $T=7384000 4504000 0 0 $X=7384000 $Y=4504000
X4301 24 4243 nand04 $T=7456000 13088000 0 0 $X=7456000 $Y=13088000
X4302 24 4244 nand04 $T=7472000 1024000 0 0 $X=7472000 $Y=1024000
X4303 24 4245 nand04 $T=7560000 2880000 0 0 $X=7560000 $Y=2880000
X4304 24 4246 nand04 $T=7592000 7984000 0 0 $X=7592000 $Y=7984000
X4305 24 4247 nand04 $T=7592000 8912000 0 0 $X=7592000 $Y=8912000
X4306 24 4248 nand04 $T=7624000 5664000 0 0 $X=7624000 $Y=5664000
X4307 24 4249 nand04 $T=7704000 11696000 0 0 $X=7704000 $Y=11696000
X4308 24 4250 nand04 $T=7785000 5664000 1 180 $X=7736000 $Y=5664000
X4309 24 4251 nand04 $T=7808000 10304000 0 0 $X=7808000 $Y=10304000
X4310 24 4252 nand04 $T=7856000 3112000 0 0 $X=7856000 $Y=3112000
X4311 24 4253 nand04 $T=8049000 1952000 1 180 $X=8000000 $Y=1952000
X4312 24 4254 nand04 $T=8057000 7752000 1 180 $X=8008000 $Y=7752000
X4313 24 4255 nand04 $T=8016000 7520000 0 0 $X=8016000 $Y=7520000
X4314 24 4256 nand04 $T=8056000 1952000 0 0 $X=8056000 $Y=1952000
X4315 24 4257 nand04 $T=8080000 2880000 0 0 $X=8080000 $Y=2880000
X4316 24 4258 nand04 $T=8128000 12392000 0 0 $X=8128000 $Y=12392000
X4317 24 4259 nand04 $T=8144000 11696000 0 0 $X=8144000 $Y=11696000
X4318 24 4260 nand04 $T=8201000 5664000 1 180 $X=8152000 $Y=5664000
X4319 24 4261 nand04 $T=8224000 1952000 0 0 $X=8224000 $Y=1952000
X4320 24 4262 nand04 $T=8240000 12392000 0 0 $X=8240000 $Y=12392000
X4321 24 4263 nand04 $T=8297000 792000 1 180 $X=8248000 $Y=792000
X4322 24 4264 nand04 $T=8297000 3808000 1 180 $X=8248000 $Y=3808000
X4323 24 4265 nand04 $T=8321000 9840000 1 180 $X=8272000 $Y=9840000
X4324 24 4266 nand04 $T=8345000 2880000 1 180 $X=8296000 $Y=2880000
X4325 24 4267 nand04 $T=8336000 10768000 0 0 $X=8336000 $Y=10768000
X4326 24 4268 nand04 $T=8360000 792000 0 0 $X=8360000 $Y=792000
X4327 24 4269 nand04 $T=8449000 9376000 1 180 $X=8400000 $Y=9376000
X4328 24 4270 nand04 $T=8416000 1024000 0 0 $X=8416000 $Y=1024000
X4329 24 4271 nand04 $T=8424000 6360000 0 0 $X=8424000 $Y=6360000
X4330 24 4272 nand04 $T=8448000 328000 0 0 $X=8448000 $Y=328000
X4331 24 4273 nand04 $T=8480000 4968000 0 0 $X=8480000 $Y=4968000
X4332 24 4274 nand04 $T=8745000 13320000 1 180 $X=8696000 $Y=13320000
X4333 24 4275 nand04 $T=8736000 7520000 0 0 $X=8736000 $Y=7520000
X4334 24 4276 nand04 $T=8736000 10304000 0 0 $X=8736000 $Y=10304000
X4335 24 4277 nand04 $T=8784000 4736000 0 0 $X=8784000 $Y=4736000
X4336 24 4278 nand04 $T=8897000 12856000 1 180 $X=8848000 $Y=12856000
X4337 24 4279 nand04 $T=9001000 3344000 1 180 $X=8952000 $Y=3344000
X4338 24 4280 nand04 $T=9009000 12392000 1 180 $X=8960000 $Y=12392000
X4339 24 4281 nand04 $T=9000000 1024000 0 0 $X=9000000 $Y=1024000
X4340 24 4282 nand04 $T=9000000 11696000 0 0 $X=9000000 $Y=11696000
X4341 24 4283 nand04 $T=9048000 4272000 0 0 $X=9048000 $Y=4272000
X4342 24 4284 nand04 $T=9121000 12392000 1 180 $X=9072000 $Y=12392000
X4343 24 4285 nand04 $T=9088000 328000 0 0 $X=9088000 $Y=328000
X4344 24 4286 nand04 $T=9096000 10536000 0 0 $X=9096000 $Y=10536000
X4345 24 4287 nand04 $T=9169000 8912000 1 180 $X=9120000 $Y=8912000
X4346 24 4288 nand04 $T=9120000 9840000 0 0 $X=9120000 $Y=9840000
X4347 24 4289 nand04 $T=9144000 6360000 0 0 $X=9144000 $Y=6360000
X4348 24 4290 nand04 $T=9200000 3808000 0 0 $X=9200000 $Y=3808000
X4349 24 4291 nand04 $T=9200000 5432000 0 0 $X=9200000 $Y=5432000
X4350 24 4292 nand04 $T=9369000 7288000 1 180 $X=9320000 $Y=7288000
X4351 24 4293 nand04 $T=9400000 1952000 0 0 $X=9400000 $Y=1952000
X4352 24 4294 nand04 $T=9457000 4040000 1 180 $X=9408000 $Y=4040000
X4353 24 4295 nand04 $T=9465000 8216000 1 180 $X=9416000 $Y=8216000
X4354 24 4296 nand04 $T=9480000 792000 0 0 $X=9480000 $Y=792000
X4355 24 4297 nand04 $T=9737000 4040000 1 180 $X=9688000 $Y=4040000
X4356 24 4298 nand04 $T=9720000 7984000 0 0 $X=9720000 $Y=7984000
X4357 24 4299 nand04 $T=9752000 1720000 0 0 $X=9752000 $Y=1720000
X4358 24 4300 nand04 $T=9792000 6128000 0 0 $X=9792000 $Y=6128000
X4359 24 2350 nand04 $T=9993000 10536000 1 180 $X=9944000 $Y=10536000
X4360 24 4301 nand04 $T=10016000 10304000 0 0 $X=10016000 $Y=10304000
X4361 24 4302 nand04 $T=10032000 1024000 0 0 $X=10032000 $Y=1024000
X4362 24 4303 nand04 $T=10048000 9376000 0 0 $X=10048000 $Y=9376000
X4363 24 4304 nand04 $T=10105000 5896000 1 180 $X=10056000 $Y=5896000
X4364 24 4305 nand04 $T=10112000 6360000 0 0 $X=10112000 $Y=6360000
X4365 24 4306 nand04 $T=10128000 9840000 0 0 $X=10128000 $Y=9840000
X4366 24 4307 nand04 $T=10201000 9144000 1 180 $X=10152000 $Y=9144000
X4367 24 4308 nand04 $T=10192000 11928000 0 0 $X=10192000 $Y=11928000
X4368 24 4309 nand04 $T=10369000 12392000 1 180 $X=10320000 $Y=12392000
X4369 24 4310 nand04 $T=10360000 1952000 0 0 $X=10360000 $Y=1952000
X4370 24 4311 nand04 $T=10360000 4504000 0 0 $X=10360000 $Y=4504000
X4371 24 4312 nand04 $T=10505000 9376000 1 180 $X=10456000 $Y=9376000
X4372 24 4313 nand04 $T=10464000 3808000 0 0 $X=10464000 $Y=3808000
X4373 24 4314 nand04 $T=10537000 7056000 1 180 $X=10488000 $Y=7056000
X4374 24 4315 nand04 $T=10520000 3808000 0 0 $X=10520000 $Y=3808000
X4375 24 4316 nand04 $T=10528000 3576000 0 0 $X=10528000 $Y=3576000
X4376 24 4317 nand04 $T=10633000 8912000 1 180 $X=10584000 $Y=8912000
X4377 24 4318 nand04 $T=10632000 7288000 0 0 $X=10632000 $Y=7288000
X4378 24 4319 nand04 $T=10737000 8216000 1 180 $X=10688000 $Y=8216000
X4379 24 4320 nand04 $T=10769000 6824000 1 180 $X=10720000 $Y=6824000
X4380 24 4321 nand04 $T=10769000 13320000 1 180 $X=10720000 $Y=13320000
X4381 24 4322 nand04 $T=10752000 5896000 0 0 $X=10752000 $Y=5896000
X4382 24 4323 nand04 $T=10809000 5200000 1 180 $X=10760000 $Y=5200000
X4383 24 4324 nand04 $T=10825000 4504000 1 180 $X=10776000 $Y=4504000
X4384 24 4325 nand04 $T=10833000 13088000 1 180 $X=10784000 $Y=13088000
X4385 24 4326 nand04 $T=10849000 6128000 1 180 $X=10800000 $Y=6128000
X4386 24 4327 nand04 $T=10824000 2184000 0 0 $X=10824000 $Y=2184000
X4387 24 4328 nand04 $T=10873000 5664000 1 180 $X=10824000 $Y=5664000
X4388 24 4329 nand04 $T=10881000 6824000 1 180 $X=10832000 $Y=6824000
X4389 24 4330 nand04 $T=10881000 11000000 1 180 $X=10832000 $Y=11000000
X4390 24 4331 nand04 $T=10913000 8216000 1 180 $X=10864000 $Y=8216000
X4391 24 4332 nand04 $T=10936000 7520000 0 0 $X=10936000 $Y=7520000
X4392 24 4333 nand04 $T=11200000 10536000 0 0 $X=11200000 $Y=10536000
X4393 24 4334 nand04 $T=11248000 6360000 0 0 $X=11248000 $Y=6360000
X4394 24 4335 nand04 $T=11345000 9144000 1 180 $X=11296000 $Y=9144000
X4395 24 4336 nand04 $T=11384000 4736000 0 0 $X=11384000 $Y=4736000
X4396 24 4337 nand04 $T=11416000 7752000 0 0 $X=11416000 $Y=7752000
X4397 24 4338 nand04 $T=11489000 9840000 1 180 $X=11440000 $Y=9840000
X4398 24 4339 nand04 $T=11537000 12624000 1 180 $X=11488000 $Y=12624000
X4399 24 4340 nand04 $T=11496000 3576000 0 0 $X=11496000 $Y=3576000
X4400 24 4341 nand04 $T=11545000 11000000 1 180 $X=11496000 $Y=11000000
X4401 24 4342 nand04 $T=11625000 2416000 1 180 $X=11576000 $Y=2416000
X4402 24 4343 nand04 $T=11625000 12392000 1 180 $X=11576000 $Y=12392000
X4403 24 4344 nand04 $T=11584000 7752000 0 0 $X=11584000 $Y=7752000
X4404 24 4345 nand04 $T=11584000 11696000 0 0 $X=11584000 $Y=11696000
X4405 24 4346 nand04 $T=11632000 2416000 0 0 $X=11632000 $Y=2416000
X4406 24 4347 nand04 $T=11744000 6592000 0 0 $X=11744000 $Y=6592000
X4407 24 4348 nand04 $T=12009000 11232000 1 180 $X=11960000 $Y=11232000
X4408 24 4349 nand04 $T=12033000 3808000 1 180 $X=11984000 $Y=3808000
X4409 24 4350 nand04 $T=12160000 4272000 0 0 $X=12160000 $Y=4272000
X4410 24 oai221 $T=10632000 1488000 0 0 $X=10632000 $Y=1488000
X4411 24 oai221 $T=11289500 1488000 1 180 $X=11224000 $Y=1488000
X4412 24 oai221 $T=11625500 1488000 1 180 $X=11560000 $Y=1488000
X4413 24 oai221 $T=11696000 560000 0 0 $X=11696000 $Y=560000
X4414 24 oai221 $T=11888000 7056000 0 0 $X=11888000 $Y=7056000
X4415 24 oai221 $T=11896000 7288000 0 0 $X=11896000 $Y=7288000
X4416 24 oai221 $T=12064000 1488000 0 0 $X=12064000 $Y=1488000
X4417 24 oai221 $T=12201500 1488000 1 180 $X=12136000 $Y=1488000
X4418 24 ICV_5 $T=5808000 12160000 1 180 $X=5624000 $Y=12160000
X4419 24 ICV_5 $T=6208000 8680000 1 180 $X=6024000 $Y=8680000
X4420 24 ICV_5 $T=6216000 4736000 1 180 $X=6032000 $Y=4736000
X4421 24 ICV_5 $T=6320000 2184000 1 180 $X=6136000 $Y=2184000
X4422 24 ICV_5 $T=6632000 5432000 1 180 $X=6448000 $Y=5432000
X4423 24 ICV_5 $T=7680000 4504000 1 180 $X=7496000 $Y=4504000
X4424 24 ICV_5 $T=9304000 4504000 1 180 $X=9120000 $Y=4504000
X4425 24 ICV_5 $T=10648000 12160000 1 180 $X=10464000 $Y=12160000
X4426 24 ICV_5 $T=11480000 13552000 1 180 $X=11296000 $Y=13552000
X4427 24 ICV_5 $T=12280000 5432000 1 180 $X=12096000 $Y=5432000
X4428 24 ICV_5 $T=12280000 8216000 1 180 $X=12096000 $Y=8216000
X4429 24 ICV_5 $T=12280000 10536000 1 180 $X=12096000 $Y=10536000
X4430 24 ICV_5 $T=12280000 11464000 1 180 $X=12096000 $Y=11464000
X4431 24 ICV_5 $T=12280000 12856000 1 180 $X=12096000 $Y=12856000
X4432 24 4351 ICV_6 $T=400000 4968000 0 0 $X=400000 $Y=4968000
X4433 24 4352 ICV_6 $T=1408000 5200000 0 0 $X=1408000 $Y=5200000
X4434 24 4353 ICV_6 $T=1568000 6360000 0 0 $X=1568000 $Y=6360000
X4435 24 4354 ICV_6 $T=1616000 4040000 0 0 $X=1616000 $Y=4040000
X4436 24 4355 ICV_6 $T=1640000 3808000 0 0 $X=1640000 $Y=3808000
X4437 24 4356 ICV_6 $T=1656000 6592000 0 0 $X=1656000 $Y=6592000
X4438 24 4357 ICV_6 $T=1664000 3576000 0 0 $X=1664000 $Y=3576000
X4439 24 4358 ICV_6 $T=1672000 5896000 0 0 $X=1672000 $Y=5896000
X4440 24 4359 ICV_6 $T=1720000 5664000 0 0 $X=1720000 $Y=5664000
X4441 24 4360 ICV_6 $T=1976000 8216000 0 0 $X=1976000 $Y=8216000
X4442 24 4361 ICV_6 $T=1992000 8448000 0 0 $X=1992000 $Y=8448000
X4443 24 4362 ICV_6 $T=2200000 6360000 0 0 $X=2200000 $Y=6360000
X4444 24 4363 ICV_6 $T=2376000 5432000 0 0 $X=2376000 $Y=5432000
X4445 24 4364 ICV_6 $T=2496000 10536000 0 0 $X=2496000 $Y=10536000
X4446 24 4365 ICV_6 $T=2712000 12160000 0 0 $X=2712000 $Y=12160000
X4447 24 4366 ICV_6 $T=2744000 10536000 0 0 $X=2744000 $Y=10536000
X4448 24 4367 ICV_6 $T=2992000 10536000 0 0 $X=2992000 $Y=10536000
X4449 24 2311 ICV_6 $T=3000000 5664000 0 0 $X=3000000 $Y=5664000
X4450 24 4368 ICV_6 $T=3056000 4504000 0 0 $X=3056000 $Y=4504000
X4451 24 4369 ICV_6 $T=3056000 4736000 0 0 $X=3056000 $Y=4736000
X4452 24 4370 ICV_6 $T=3064000 3112000 0 0 $X=3064000 $Y=3112000
X4453 24 4371 ICV_6 $T=3144000 1024000 0 0 $X=3144000 $Y=1024000
X4454 24 4372 ICV_6 $T=3152000 3344000 0 0 $X=3152000 $Y=3344000
X4455 24 4373 ICV_6 $T=3152000 9376000 0 0 $X=3152000 $Y=9376000
X4456 24 4374 ICV_6 $T=3192000 6360000 0 0 $X=3192000 $Y=6360000
X4457 24 4375 ICV_6 $T=3200000 560000 0 0 $X=3200000 $Y=560000
X4458 24 4376 ICV_6 $T=3240000 10536000 0 0 $X=3240000 $Y=10536000
X4459 24 4377 ICV_6 $T=3248000 5664000 0 0 $X=3248000 $Y=5664000
X4460 24 4378 ICV_6 $T=3248000 8912000 0 0 $X=3248000 $Y=8912000
X4461 24 4379 ICV_6 $T=3280000 792000 0 0 $X=3280000 $Y=792000
X4462 24 4380 ICV_6 $T=3312000 5896000 0 0 $X=3312000 $Y=5896000
X4463 24 4381 ICV_6 $T=3384000 1256000 0 0 $X=3384000 $Y=1256000
X4464 24 4382 ICV_6 $T=3400000 3344000 0 0 $X=3400000 $Y=3344000
X4465 24 4383 ICV_6 $T=3432000 1720000 0 0 $X=3432000 $Y=1720000
X4466 24 4384 ICV_6 $T=3448000 560000 0 0 $X=3448000 $Y=560000
X4467 24 4385 ICV_6 $T=3456000 1024000 0 0 $X=3456000 $Y=1024000
X4468 24 4386 ICV_6 $T=3488000 10536000 0 0 $X=3488000 $Y=10536000
X4469 24 4387 ICV_6 $T=3512000 2184000 0 0 $X=3512000 $Y=2184000
X4470 24 4388 ICV_6 $T=3632000 1256000 0 0 $X=3632000 $Y=1256000
X4471 24 4389 ICV_6 $T=3840000 8448000 0 0 $X=3840000 $Y=8448000
X4472 24 4390 ICV_6 $T=4200000 1952000 0 0 $X=4200000 $Y=1952000
X4473 24 4391 ICV_6 $T=4208000 2880000 0 0 $X=4208000 $Y=2880000
X4474 24 4392 ICV_6 $T=4248000 1488000 0 0 $X=4248000 $Y=1488000
X4475 24 4393 ICV_6 $T=4384000 4272000 0 0 $X=4384000 $Y=4272000
X4476 24 4394 ICV_6 $T=4400000 8448000 0 0 $X=4400000 $Y=8448000
X4477 24 4395 ICV_6 $T=4432000 3344000 0 0 $X=4432000 $Y=3344000
X4478 24 4396 ICV_6 $T=4448000 3808000 0 0 $X=4448000 $Y=3808000
X4479 24 4397 ICV_6 $T=4456000 2880000 0 0 $X=4456000 $Y=2880000
X4480 24 4398 ICV_6 $T=4496000 3576000 0 0 $X=4496000 $Y=3576000
X4481 24 4399 ICV_6 $T=4528000 6824000 0 0 $X=4528000 $Y=6824000
X4482 24 4400 ICV_6 $T=4552000 3112000 0 0 $X=4552000 $Y=3112000
X4483 24 4401 ICV_6 $T=4560000 9608000 0 0 $X=4560000 $Y=9608000
X4484 24 4402 ICV_6 $T=4584000 96000 0 0 $X=4584000 $Y=96000
X4485 24 4403 ICV_6 $T=4584000 2416000 0 0 $X=4584000 $Y=2416000
X4486 24 4404 ICV_6 $T=4632000 4272000 0 0 $X=4632000 $Y=4272000
X4487 24 4405 ICV_6 $T=4648000 8448000 0 0 $X=4648000 $Y=8448000
X4488 24 4406 ICV_6 $T=4696000 3808000 0 0 $X=4696000 $Y=3808000
X4489 24 4407 ICV_6 $T=4704000 2880000 0 0 $X=4704000 $Y=2880000
X4490 24 4408 ICV_6 $T=4800000 7288000 0 0 $X=4800000 $Y=7288000
X4491 24 4409 ICV_6 $T=4816000 2648000 0 0 $X=4816000 $Y=2648000
X4492 24 4410 ICV_6 $T=4840000 328000 0 0 $X=4840000 $Y=328000
X4493 24 4411 ICV_6 $T=4848000 4040000 0 0 $X=4848000 $Y=4040000
X4494 24 4412 ICV_6 $T=4872000 1488000 0 0 $X=4872000 $Y=1488000
X4495 24 4413 ICV_6 $T=4880000 2184000 0 0 $X=4880000 $Y=2184000
X4496 24 4414 ICV_6 $T=4984000 1952000 0 0 $X=4984000 $Y=1952000
X4497 24 4415 ICV_6 $T=5048000 7288000 0 0 $X=5048000 $Y=7288000
X4498 24 4416 ICV_6 $T=5056000 7056000 0 0 $X=5056000 $Y=7056000
X4499 24 4417 ICV_6 $T=5120000 1488000 0 0 $X=5120000 $Y=1488000
X4500 24 4418 ICV_6 $T=5128000 2184000 0 0 $X=5128000 $Y=2184000
X4501 24 4419 ICV_6 $T=5136000 7520000 0 0 $X=5136000 $Y=7520000
X4502 24 4420 ICV_6 $T=5304000 11696000 0 0 $X=5304000 $Y=11696000
X4503 24 4421 ICV_6 $T=5368000 1488000 0 0 $X=5368000 $Y=1488000
X4504 24 4422 ICV_6 $T=5440000 1720000 0 0 $X=5440000 $Y=1720000
X4505 24 4423 ICV_6 $T=5480000 8216000 0 0 $X=5480000 $Y=8216000
X4506 24 4424 ICV_6 $T=5512000 1952000 0 0 $X=5512000 $Y=1952000
X4507 24 4425 ICV_6 $T=5552000 1256000 0 0 $X=5552000 $Y=1256000
X4508 24 4426 ICV_6 $T=5616000 1488000 0 0 $X=5616000 $Y=1488000
X4509 24 4427 ICV_6 $T=5824000 2184000 0 0 $X=5824000 $Y=2184000
X4510 24 4428 ICV_6 $T=5864000 1488000 0 0 $X=5864000 $Y=1488000
X4511 24 4429 ICV_6 $T=5904000 7520000 0 0 $X=5904000 $Y=7520000
X4512 24 4430 ICV_6 $T=5936000 328000 0 0 $X=5936000 $Y=328000
X4513 24 4431 ICV_6 $T=6104000 1256000 0 0 $X=6104000 $Y=1256000
X4514 24 4432 ICV_6 $T=6128000 7288000 0 0 $X=6128000 $Y=7288000
X4515 24 4433 ICV_6 $T=6224000 10536000 0 0 $X=6224000 $Y=10536000
X4516 24 4434 ICV_6 $T=6248000 4968000 0 0 $X=6248000 $Y=4968000
X4517 24 4435 ICV_6 $T=6320000 3808000 0 0 $X=6320000 $Y=3808000
X4518 24 4436 ICV_6 $T=6320000 13552000 0 0 $X=6320000 $Y=13552000
X4519 24 4437 ICV_6 $T=6328000 4040000 0 0 $X=6328000 $Y=4040000
X4520 24 4438 ICV_6 $T=6352000 1256000 0 0 $X=6352000 $Y=1256000
X4521 24 4439 ICV_6 $T=6360000 11464000 0 0 $X=6360000 $Y=11464000
X4522 24 4440 ICV_6 $T=6376000 7288000 0 0 $X=6376000 $Y=7288000
X4523 24 4441 ICV_6 $T=6400000 11696000 0 0 $X=6400000 $Y=11696000
X4524 24 4442 ICV_6 $T=6408000 11000000 0 0 $X=6408000 $Y=11000000
X4525 24 4443 ICV_6 $T=6424000 1488000 0 0 $X=6424000 $Y=1488000
X4526 24 4444 ICV_6 $T=6424000 4272000 0 0 $X=6424000 $Y=4272000
X4527 24 4445 ICV_6 $T=6432000 7984000 0 0 $X=6432000 $Y=7984000
X4528 24 4446 ICV_6 $T=6456000 9608000 0 0 $X=6456000 $Y=9608000
X4529 24 4447 ICV_6 $T=6472000 10536000 0 0 $X=6472000 $Y=10536000
X4530 24 4448 ICV_6 $T=6480000 792000 0 0 $X=6480000 $Y=792000
X4531 24 4449 ICV_6 $T=6504000 12624000 0 0 $X=6504000 $Y=12624000
X4532 24 4450 ICV_6 $T=6568000 3808000 0 0 $X=6568000 $Y=3808000
X4533 24 4451 ICV_6 $T=6576000 4040000 0 0 $X=6576000 $Y=4040000
X4534 24 4452 ICV_6 $T=6584000 7520000 0 0 $X=6584000 $Y=7520000
X4535 24 4453 ICV_6 $T=6584000 7752000 0 0 $X=6584000 $Y=7752000
X4536 24 4454 ICV_6 $T=6624000 7288000 0 0 $X=6624000 $Y=7288000
X4537 24 4455 ICV_6 $T=6640000 5200000 0 0 $X=6640000 $Y=5200000
X4538 24 4456 ICV_6 $T=6728000 560000 0 0 $X=6728000 $Y=560000
X4539 24 4457 ICV_6 $T=6752000 12624000 0 0 $X=6752000 $Y=12624000
X4540 24 4458 ICV_6 $T=6808000 13552000 0 0 $X=6808000 $Y=13552000
X4541 24 4459 ICV_6 $T=6824000 4040000 0 0 $X=6824000 $Y=4040000
X4542 24 4460 ICV_6 $T=6832000 1720000 0 0 $X=6832000 $Y=1720000
X4543 24 4461 ICV_6 $T=6840000 1952000 0 0 $X=6840000 $Y=1952000
X4544 24 4462 ICV_6 $T=6848000 8448000 0 0 $X=6848000 $Y=8448000
X4545 24 4463 ICV_6 $T=6864000 2416000 0 0 $X=6864000 $Y=2416000
X4546 24 4464 ICV_6 $T=6888000 5200000 0 0 $X=6888000 $Y=5200000
X4547 24 4465 ICV_6 $T=6896000 5664000 0 0 $X=6896000 $Y=5664000
X4548 24 4466 ICV_6 $T=7008000 5432000 0 0 $X=7008000 $Y=5432000
X4549 24 4467 ICV_6 $T=7120000 13552000 0 0 $X=7120000 $Y=13552000
X4550 24 4468 ICV_6 $T=7136000 5200000 0 0 $X=7136000 $Y=5200000
X4551 24 4469 ICV_6 $T=7200000 10536000 0 0 $X=7200000 $Y=10536000
X4552 24 4470 ICV_6 $T=7224000 3576000 0 0 $X=7224000 $Y=3576000
X4553 24 4471 ICV_6 $T=7312000 6592000 0 0 $X=7312000 $Y=6592000
X4554 24 4472 ICV_6 $T=7344000 560000 0 0 $X=7344000 $Y=560000
X4555 24 4473 ICV_6 $T=7352000 6360000 0 0 $X=7352000 $Y=6360000
X4556 24 4474 ICV_6 $T=7384000 5200000 0 0 $X=7384000 $Y=5200000
X4557 24 4475 ICV_6 $T=7416000 10768000 0 0 $X=7416000 $Y=10768000
X4558 24 4476 ICV_6 $T=7560000 6592000 0 0 $X=7560000 $Y=6592000
X4559 24 4477 ICV_6 $T=7568000 1720000 0 0 $X=7568000 $Y=1720000
X4560 24 4478 ICV_6 $T=7584000 792000 0 0 $X=7584000 $Y=792000
X4561 24 4479 ICV_6 $T=7600000 6360000 0 0 $X=7600000 $Y=6360000
X4562 24 4480 ICV_6 $T=7656000 4736000 0 0 $X=7656000 $Y=4736000
X4563 24 4481 ICV_6 $T=7680000 328000 0 0 $X=7680000 $Y=328000
X4564 24 4482 ICV_6 $T=7744000 96000 0 0 $X=7744000 $Y=96000
X4565 24 4483 ICV_6 $T=7744000 4504000 0 0 $X=7744000 $Y=4504000
X4566 24 4484 ICV_6 $T=7808000 6592000 0 0 $X=7808000 $Y=6592000
X4567 24 4485 ICV_6 $T=7928000 328000 0 0 $X=7928000 $Y=328000
X4568 24 4486 ICV_6 $T=7944000 1256000 0 0 $X=7944000 $Y=1256000
X4569 24 4487 ICV_6 $T=7944000 5432000 0 0 $X=7944000 $Y=5432000
X4570 24 4488 ICV_6 $T=7992000 96000 0 0 $X=7992000 $Y=96000
X4571 24 4489 ICV_6 $T=7992000 4504000 0 0 $X=7992000 $Y=4504000
X4572 24 4490 ICV_6 $T=8168000 1024000 0 0 $X=8168000 $Y=1024000
X4573 24 4491 ICV_6 $T=8240000 96000 0 0 $X=8240000 $Y=96000
X4574 24 4492 ICV_6 $T=8304000 11464000 0 0 $X=8304000 $Y=11464000
X4575 24 4493 ICV_6 $T=8360000 6592000 0 0 $X=8360000 $Y=6592000
X4576 24 4494 ICV_6 $T=8424000 10768000 0 0 $X=8424000 $Y=10768000
X4577 24 4495 ICV_6 $T=8440000 6128000 0 0 $X=8440000 $Y=6128000
X4578 24 4496 ICV_6 $T=8560000 4272000 0 0 $X=8560000 $Y=4272000
X4579 24 4497 ICV_6 $T=8608000 5200000 0 0 $X=8608000 $Y=5200000
X4580 24 4498 ICV_6 $T=8624000 5432000 0 0 $X=8624000 $Y=5432000
X4581 24 4499 ICV_6 $T=8672000 10768000 0 0 $X=8672000 $Y=10768000
X4582 24 4500 ICV_6 $T=8768000 96000 0 0 $X=8768000 $Y=96000
X4583 24 4501 ICV_6 $T=8776000 4968000 0 0 $X=8776000 $Y=4968000
X4584 24 4502 ICV_6 $T=8776000 9608000 0 0 $X=8776000 $Y=9608000
X4585 24 4503 ICV_6 $T=8816000 11000000 0 0 $X=8816000 $Y=11000000
X4586 24 4504 ICV_6 $T=8856000 5200000 0 0 $X=8856000 $Y=5200000
X4587 24 4505 ICV_6 $T=8960000 4736000 0 0 $X=8960000 $Y=4736000
X4588 24 4506 ICV_6 $T=9024000 4968000 0 0 $X=9024000 $Y=4968000
X4589 24 4507 ICV_6 $T=9024000 9608000 0 0 $X=9024000 $Y=9608000
X4590 24 4508 ICV_6 $T=9040000 6592000 0 0 $X=9040000 $Y=6592000
X4591 24 4509 ICV_6 $T=9120000 11696000 0 0 $X=9120000 $Y=11696000
X4592 24 4510 ICV_6 $T=9288000 6592000 0 0 $X=9288000 $Y=6592000
X4593 24 4511 ICV_6 $T=9296000 1488000 0 0 $X=9296000 $Y=1488000
X4594 24 4512 ICV_6 $T=9296000 2880000 0 0 $X=9296000 $Y=2880000
X4595 24 4513 ICV_6 $T=9320000 6360000 0 0 $X=9320000 $Y=6360000
X4596 24 4514 ICV_6 $T=9328000 5896000 0 0 $X=9328000 $Y=5896000
X4597 24 4515 ICV_6 $T=9536000 1256000 0 0 $X=9536000 $Y=1256000
X4598 24 4516 ICV_6 $T=9568000 6360000 0 0 $X=9568000 $Y=6360000
X4599 24 4517 ICV_6 $T=9648000 7520000 0 0 $X=9648000 $Y=7520000
X4600 24 4518 ICV_6 $T=9760000 4736000 0 0 $X=9760000 $Y=4736000
X4601 24 4519 ICV_6 $T=9808000 1720000 0 0 $X=9808000 $Y=1720000
X4602 24 4520 ICV_6 $T=9848000 1488000 0 0 $X=9848000 $Y=1488000
X4603 24 4521 ICV_6 $T=9872000 328000 0 0 $X=9872000 $Y=328000
X4604 24 4522 ICV_6 $T=9880000 2648000 0 0 $X=9880000 $Y=2648000
X4605 24 4523 ICV_6 $T=9888000 6592000 0 0 $X=9888000 $Y=6592000
X4606 24 4524 ICV_6 $T=9904000 2416000 0 0 $X=9904000 $Y=2416000
X4607 24 4525 ICV_6 $T=9928000 3808000 0 0 $X=9928000 $Y=3808000
X4608 24 4526 ICV_6 $T=9952000 6824000 0 0 $X=9952000 $Y=6824000
X4609 24 4527 ICV_6 $T=9960000 10768000 0 0 $X=9960000 $Y=10768000
X4610 24 4528 ICV_6 $T=9992000 3576000 0 0 $X=9992000 $Y=3576000
X4611 24 4529 ICV_6 $T=10000000 7056000 0 0 $X=10000000 $Y=7056000
X4612 24 4530 ICV_6 $T=10040000 3112000 0 0 $X=10040000 $Y=3112000
X4613 24 4531 ICV_6 $T=10104000 4968000 0 0 $X=10104000 $Y=4968000
X4614 24 4532 ICV_6 $T=10184000 10304000 0 0 $X=10184000 $Y=10304000
X4615 24 4533 ICV_6 $T=10248000 2416000 0 0 $X=10248000 $Y=2416000
X4616 24 4534 ICV_6 $T=10344000 13552000 0 0 $X=10344000 $Y=13552000
X4617 24 4535 ICV_6 $T=10424000 10536000 0 0 $X=10424000 $Y=10536000
X4618 24 4536 ICV_6 $T=10424000 11928000 0 0 $X=10424000 $Y=11928000
X4619 24 4537 ICV_6 $T=10496000 2416000 0 0 $X=10496000 $Y=2416000
X4620 24 4538 ICV_6 $T=10496000 12392000 0 0 $X=10496000 $Y=12392000
X4621 24 4539 ICV_6 $T=10536000 8680000 0 0 $X=10536000 $Y=8680000
X4622 24 4540 ICV_6 $T=10640000 3344000 0 0 $X=10640000 $Y=3344000
X4623 24 4541 ICV_6 $T=10640000 12624000 0 0 $X=10640000 $Y=12624000
X4624 24 4542 ICV_6 $T=10656000 4968000 0 0 $X=10656000 $Y=4968000
X4625 24 4543 ICV_6 $T=10712000 12160000 0 0 $X=10712000 $Y=12160000
X4626 24 4544 ICV_6 $T=10824000 3576000 0 0 $X=10824000 $Y=3576000
X4627 24 4545 ICV_6 $T=10936000 5200000 0 0 $X=10936000 $Y=5200000
X4628 24 4546 ICV_6 $T=11040000 2648000 0 0 $X=11040000 $Y=2648000
X4629 24 4102 ICV_6 $T=11040000 11928000 0 0 $X=11040000 $Y=11928000
X4630 24 4547 ICV_6 $T=11056000 7288000 0 0 $X=11056000 $Y=7288000
X4631 24 4548 ICV_6 $T=11056000 7520000 0 0 $X=11056000 $Y=7520000
X4632 24 4549 ICV_6 $T=11088000 8680000 0 0 $X=11088000 $Y=8680000
X4633 24 4550 ICV_6 $T=11112000 2880000 0 0 $X=11112000 $Y=2880000
X4634 24 4551 ICV_6 $T=11280000 7056000 0 0 $X=11280000 $Y=7056000
X4635 24 4552 ICV_6 $T=11288000 11928000 0 0 $X=11288000 $Y=11928000
X4636 24 4553 ICV_6 $T=11304000 4272000 0 0 $X=11304000 $Y=4272000
X4637 24 4554 ICV_6 $T=11304000 7520000 0 0 $X=11304000 $Y=7520000
X4638 24 4555 ICV_6 $T=11320000 6128000 0 0 $X=11320000 $Y=6128000
X4639 24 4556 ICV_6 $T=11400000 4968000 0 0 $X=11400000 $Y=4968000
X4640 24 4557 ICV_6 $T=11536000 11928000 0 0 $X=11536000 $Y=11928000
X4641 24 4558 ICV_6 $T=11552000 11464000 0 0 $X=11552000 $Y=11464000
X4642 24 4559 ICV_6 $T=11568000 6128000 0 0 $X=11568000 $Y=6128000
X4643 24 4560 ICV_6 $T=11592000 9608000 0 0 $X=11592000 $Y=9608000
X4644 24 4561 ICV_6 $T=11600000 5200000 0 0 $X=11600000 $Y=5200000
X4645 24 4562 ICV_6 $T=11608000 7288000 0 0 $X=11608000 $Y=7288000
X4646 24 4563 ICV_6 $T=11736000 4736000 0 0 $X=11736000 $Y=4736000
X4647 24 4564 ICV_6 $T=11784000 2648000 0 0 $X=11784000 $Y=2648000
X4648 24 4565 ICV_6 $T=11792000 4968000 0 0 $X=11792000 $Y=4968000
X4649 24 4566 ICV_6 $T=11792000 12392000 0 0 $X=11792000 $Y=12392000
X4650 24 4567 ICV_6 $T=11848000 2880000 0 0 $X=11848000 $Y=2880000
X4651 24 4568 ICV_6 $T=11848000 4040000 0 0 $X=11848000 $Y=4040000
X4652 24 4569 ICV_6 $T=11912000 4504000 0 0 $X=11912000 $Y=4504000
X4653 24 4570 ICV_6 $T=12032000 2648000 0 0 $X=12032000 $Y=2648000
X4654 24 4571 ICV_6 $T=12096000 2184000 0 0 $X=12096000 $Y=2184000
X4655 24 4572 ICV_6 $T=12096000 2416000 0 0 $X=12096000 $Y=2416000
X4656 24 4573 ICV_6 $T=12096000 3112000 0 0 $X=12096000 $Y=3112000
X4657 24 4574 ICV_6 $T=12096000 11696000 0 0 $X=12096000 $Y=11696000
X4658 24 4575 ICV_7 $T=336000 5200000 1 180 $X=152000 $Y=5200000
X4659 24 3682 ICV_7 $T=888000 5896000 1 180 $X=704000 $Y=5896000
X4660 24 3922 ICV_7 $T=7272000 6128000 1 180 $X=7088000 $Y=6128000
X4661 24 4576 ICV_7 $T=8808000 5664000 1 180 $X=8624000 $Y=5664000
X4662 24 4577 ICV_7 $T=11184000 1952000 1 180 $X=11000000 $Y=1952000
X4663 24 4578 ICV_7 $T=12280000 4040000 1 180 $X=12096000 $Y=4040000
X4664 24 ICV_8 $T=152000 8680000 0 0 $X=152000 $Y=8680000
X4665 24 ICV_8 $T=192000 9608000 0 0 $X=192000 $Y=9608000
X4666 24 ICV_8 $T=296000 9840000 0 0 $X=296000 $Y=9840000
X4667 24 ICV_8 $T=632000 13320000 0 0 $X=632000 $Y=13320000
X4668 24 ICV_8 $T=720000 9840000 0 0 $X=720000 $Y=9840000
X4669 24 ICV_8 $T=1536000 13552000 0 0 $X=1536000 $Y=13552000
X4670 24 ICV_8 $T=2664000 13088000 0 0 $X=2664000 $Y=13088000
X4671 24 ICV_8 $T=2960000 12160000 0 0 $X=2960000 $Y=12160000
X4672 24 ICV_8 $T=2968000 10768000 0 0 $X=2968000 $Y=10768000
X4673 24 ICV_8 $T=3240000 11696000 0 0 $X=3240000 $Y=11696000
X4674 24 ICV_8 $T=3472000 10304000 0 0 $X=3472000 $Y=10304000
X4675 24 ICV_8 $T=4120000 10304000 0 0 $X=4120000 $Y=10304000
X4676 24 ICV_8 $T=4920000 13320000 0 0 $X=4920000 $Y=13320000
X4677 24 ICV_8 $T=5400000 12160000 0 0 $X=5400000 $Y=12160000
X4678 24 ICV_8 $T=5696000 12856000 0 0 $X=5696000 $Y=12856000
X4679 24 ICV_8 $T=6120000 11000000 0 0 $X=6120000 $Y=11000000
X4680 24 ICV_8 $T=6192000 10768000 0 0 $X=6192000 $Y=10768000
X4681 24 ICV_8 $T=6248000 10304000 0 0 $X=6248000 $Y=10304000
X4682 24 ICV_8 $T=7328000 11000000 0 0 $X=7328000 $Y=11000000
X4683 24 ICV_8 $T=11080000 12856000 0 0 $X=11080000 $Y=12856000
X4684 24 ICV_8 $T=11544000 13552000 0 0 $X=11544000 $Y=13552000
X4685 24 ICV_8 $T=11704000 13088000 0 0 $X=11704000 $Y=13088000
X4686 24 ICV_8 $T=11912000 12624000 0 0 $X=11912000 $Y=12624000
X4687 24 ICV_8 $T=12040000 12392000 0 0 $X=12040000 $Y=12392000
X4688 24 ICV_8 $T=12056000 12160000 0 0 $X=12056000 $Y=12160000
X4689 24 4579 ICV_9 $T=680000 11696000 0 0 $X=680000 $Y=11696000
X4690 24 4580 ICV_9 $T=984000 4968000 0 0 $X=984000 $Y=4968000
X4691 24 4581 ICV_9 $T=1048000 11232000 0 0 $X=1048000 $Y=11232000
X4692 24 4582 ICV_9 $T=1048000 13088000 0 0 $X=1048000 $Y=13088000
X4693 24 4583 ICV_9 $T=1448000 11232000 0 0 $X=1448000 $Y=11232000
X4694 24 4584 ICV_9 $T=1632000 7288000 0 0 $X=1632000 $Y=7288000
X4695 24 4585 ICV_9 $T=1632000 7984000 0 0 $X=1632000 $Y=7984000
X4696 24 4586 ICV_9 $T=1688000 8448000 0 0 $X=1688000 $Y=8448000
X4697 24 4587 ICV_9 $T=1752000 7520000 0 0 $X=1752000 $Y=7520000
X4698 24 4588 ICV_9 $T=1768000 5432000 0 0 $X=1768000 $Y=5432000
X4699 24 4589 ICV_9 $T=1840000 6360000 0 0 $X=1840000 $Y=6360000
X4700 24 4590 ICV_9 $T=1896000 4968000 0 0 $X=1896000 $Y=4968000
X4701 24 4591 ICV_9 $T=1912000 3576000 0 0 $X=1912000 $Y=3576000
X4702 24 4592 ICV_9 $T=2168000 6128000 0 0 $X=2168000 $Y=6128000
X4703 24 4593 ICV_9 $T=2176000 13088000 0 0 $X=2176000 $Y=13088000
X4704 24 4594 ICV_9 $T=2352000 7752000 0 0 $X=2352000 $Y=7752000
X4705 24 4595 ICV_9 $T=2472000 4040000 0 0 $X=2472000 $Y=4040000
X4706 24 4596 ICV_9 $T=2632000 4272000 0 0 $X=2632000 $Y=4272000
X4707 24 4597 ICV_9 $T=2736000 8680000 0 0 $X=2736000 $Y=8680000
X4708 24 4598 ICV_9 $T=2816000 3344000 0 0 $X=2816000 $Y=3344000
X4709 24 4599 ICV_9 $T=3024000 13320000 0 0 $X=3024000 $Y=13320000
X4710 24 4600 ICV_9 $T=3080000 12856000 0 0 $X=3080000 $Y=12856000
X4711 24 4601 ICV_9 $T=3400000 9376000 0 0 $X=3400000 $Y=9376000
X4712 24 4602 ICV_9 $T=3544000 3808000 0 0 $X=3544000 $Y=3808000
X4713 24 4603 ICV_9 $T=3560000 5896000 0 0 $X=3560000 $Y=5896000
X4714 24 4604 ICV_9 $T=3744000 4272000 0 0 $X=3744000 $Y=4272000
X4715 24 4605 ICV_9 $T=3776000 11696000 0 0 $X=3776000 $Y=11696000
X4716 24 4606 ICV_9 $T=3784000 1952000 0 0 $X=3784000 $Y=1952000
X4717 24 4607 ICV_9 $T=3792000 6592000 0 0 $X=3792000 $Y=6592000
X4718 24 4608 ICV_9 $T=3824000 4040000 0 0 $X=3824000 $Y=4040000
X4719 24 4609 ICV_9 $T=3840000 7520000 0 0 $X=3840000 $Y=7520000
X4720 24 4610 ICV_9 $T=3848000 2416000 0 0 $X=3848000 $Y=2416000
X4721 24 4611 ICV_9 $T=3848000 3808000 0 0 $X=3848000 $Y=3808000
X4722 24 4612 ICV_9 $T=3880000 1256000 0 0 $X=3880000 $Y=1256000
X4723 24 4613 ICV_9 $T=3880000 11928000 0 0 $X=3880000 $Y=11928000
X4724 24 4614 ICV_9 $T=3912000 6824000 0 0 $X=3912000 $Y=6824000
X4725 24 4615 ICV_9 $T=4096000 7752000 0 0 $X=4096000 $Y=7752000
X4726 24 4616 ICV_9 $T=4232000 13320000 0 0 $X=4232000 $Y=13320000
X4727 24 4617 ICV_9 $T=4296000 11464000 0 0 $X=4296000 $Y=11464000
X4728 24 4618 ICV_9 $T=4448000 1952000 0 0 $X=4448000 $Y=1952000
X4729 24 4619 ICV_9 $T=4616000 13320000 0 0 $X=4616000 $Y=13320000
X4730 24 4620 ICV_9 $T=4712000 4968000 0 0 $X=4712000 $Y=4968000
X4731 24 4621 ICV_9 $T=4752000 7056000 0 0 $X=4752000 $Y=7056000
X4732 24 4622 ICV_9 $T=4808000 9608000 0 0 $X=4808000 $Y=9608000
X4733 24 4623 ICV_9 $T=4832000 7520000 0 0 $X=4832000 $Y=7520000
X4734 24 4624 ICV_9 $T=4832000 8912000 0 0 $X=4832000 $Y=8912000
X4735 24 4625 ICV_9 $T=5224000 3808000 0 0 $X=5224000 $Y=3808000
X4736 24 4626 ICV_9 $T=5272000 6824000 0 0 $X=5272000 $Y=6824000
X4737 24 4627 ICV_9 $T=5384000 7520000 0 0 $X=5384000 $Y=7520000
X4738 24 4628 ICV_9 $T=5392000 2416000 0 0 $X=5392000 $Y=2416000
X4739 24 4629 ICV_9 $T=5472000 11000000 0 0 $X=5472000 $Y=11000000
X4740 24 4630 ICV_9 $T=5728000 8216000 0 0 $X=5728000 $Y=8216000
X4741 24 4631 ICV_9 $T=5800000 1256000 0 0 $X=5800000 $Y=1256000
X4742 24 4632 ICV_9 $T=5864000 560000 0 0 $X=5864000 $Y=560000
X4743 24 4633 ICV_9 $T=5864000 9144000 0 0 $X=5864000 $Y=9144000
X4744 24 4634 ICV_9 $T=5880000 6824000 0 0 $X=5880000 $Y=6824000
X4745 24 4635 ICV_9 $T=5904000 9840000 0 0 $X=5904000 $Y=9840000
X4746 24 4636 ICV_9 $T=6080000 3344000 0 0 $X=6080000 $Y=3344000
X4747 24 4637 ICV_9 $T=6384000 2184000 0 0 $X=6384000 $Y=2184000
X4748 24 4638 ICV_9 $T=6496000 4968000 0 0 $X=6496000 $Y=4968000
X4749 24 4639 ICV_9 $T=6504000 3344000 0 0 $X=6504000 $Y=3344000
X4750 24 4640 ICV_9 $T=6648000 11696000 0 0 $X=6648000 $Y=11696000
X4751 24 4641 ICV_9 $T=6720000 96000 0 0 $X=6720000 $Y=96000
X4752 24 4642 ICV_9 $T=6816000 3808000 0 0 $X=6816000 $Y=3808000
X4753 24 4643 ICV_9 $T=6944000 328000 0 0 $X=6944000 $Y=328000
X4754 24 4644 ICV_9 $T=6976000 13088000 0 0 $X=6976000 $Y=13088000
X4755 24 4645 ICV_9 $T=7000000 12624000 0 0 $X=7000000 $Y=12624000
X4756 24 4646 ICV_9 $T=7016000 10072000 0 0 $X=7016000 $Y=10072000
X4757 24 4647 ICV_9 $T=7048000 1024000 0 0 $X=7048000 $Y=1024000
X4758 24 4648 ICV_9 $T=7088000 1952000 0 0 $X=7088000 $Y=1952000
X4759 24 4649 ICV_9 $T=7088000 3344000 0 0 $X=7088000 $Y=3344000
X4760 24 4650 ICV_9 $T=7192000 9608000 0 0 $X=7192000 $Y=9608000
X4761 24 4651 ICV_9 $T=7272000 3112000 0 0 $X=7272000 $Y=3112000
X4762 24 4652 ICV_9 $T=7352000 9840000 0 0 $X=7352000 $Y=9840000
X4763 24 4653 ICV_9 $T=7392000 1256000 0 0 $X=7392000 $Y=1256000
X4764 24 4654 ICV_9 $T=7400000 8448000 0 0 $X=7400000 $Y=8448000
X4765 24 4655 ICV_9 $T=7472000 3576000 0 0 $X=7472000 $Y=3576000
X4766 24 4656 ICV_9 $T=7544000 12160000 0 0 $X=7544000 $Y=12160000
X4767 24 4657 ICV_9 $T=7640000 8448000 0 0 $X=7640000 $Y=8448000
X4768 24 4658 ICV_9 $T=7664000 9144000 0 0 $X=7664000 $Y=9144000
X4769 24 4659 ICV_9 $T=7728000 10768000 0 0 $X=7728000 $Y=10768000
X4770 24 4660 ICV_9 $T=7832000 12856000 0 0 $X=7832000 $Y=12856000
X4771 24 4661 ICV_9 $T=8000000 11464000 0 0 $X=8000000 $Y=11464000
X4772 24 4662 ICV_9 $T=8048000 11232000 0 0 $X=8048000 $Y=11232000
X4773 24 4663 ICV_9 $T=8056000 3576000 0 0 $X=8056000 $Y=3576000
X4774 24 4664 ICV_9 $T=8128000 1488000 0 0 $X=8128000 $Y=1488000
X4775 24 4665 ICV_9 $T=8128000 6360000 0 0 $X=8128000 $Y=6360000
X4776 24 4666 ICV_9 $T=8128000 7984000 0 0 $X=8128000 $Y=7984000
X4777 24 4667 ICV_9 $T=8184000 10536000 0 0 $X=8184000 $Y=10536000
X4778 24 4668 ICV_9 $T=8192000 5432000 0 0 $X=8192000 $Y=5432000
X4779 24 4669 ICV_9 $T=8192000 7520000 0 0 $X=8192000 $Y=7520000
X4780 24 4670 ICV_9 $T=8224000 3112000 0 0 $X=8224000 $Y=3112000
X4781 24 4671 ICV_9 $T=8256000 1256000 0 0 $X=8256000 $Y=1256000
X4782 24 4672 ICV_9 $T=8376000 560000 0 0 $X=8376000 $Y=560000
X4783 24 4673 ICV_9 $T=8384000 5664000 0 0 $X=8384000 $Y=5664000
X4784 24 4674 ICV_9 $T=8432000 1488000 0 0 $X=8432000 $Y=1488000
X4785 24 4675 ICV_9 $T=8472000 8216000 0 0 $X=8472000 $Y=8216000
X4786 24 4676 ICV_9 $T=8552000 10536000 0 0 $X=8552000 $Y=10536000
X4787 24 4677 ICV_9 $T=8560000 792000 0 0 $X=8560000 $Y=792000
X4788 24 4678 ICV_9 $T=8608000 12856000 0 0 $X=8608000 $Y=12856000
X4789 24 4679 ICV_9 $T=8664000 6360000 0 0 $X=8664000 $Y=6360000
X4790 24 4680 ICV_9 $T=8856000 10304000 0 0 $X=8856000 $Y=10304000
X4791 24 4681 ICV_9 $T=8880000 9376000 0 0 $X=8880000 $Y=9376000
X4792 24 4682 ICV_9 $T=8920000 10768000 0 0 $X=8920000 $Y=10768000
X4793 24 4683 ICV_9 $T=9016000 96000 0 0 $X=9016000 $Y=96000
X4794 24 4684 ICV_9 $T=9056000 3112000 0 0 $X=9056000 $Y=3112000
X4795 24 4685 ICV_9 $T=9056000 4040000 0 0 $X=9056000 $Y=4040000
X4796 24 4686 ICV_9 $T=9064000 6128000 0 0 $X=9064000 $Y=6128000
X4797 24 4687 ICV_9 $T=9072000 3344000 0 0 $X=9072000 $Y=3344000
X4798 24 4688 ICV_9 $T=9104000 5200000 0 0 $X=9104000 $Y=5200000
X4799 24 4689 ICV_9 $T=9112000 560000 0 0 $X=9112000 $Y=560000
X4800 24 4690 ICV_9 $T=9208000 328000 0 0 $X=9208000 $Y=328000
X4801 24 4691 ICV_9 $T=9232000 7056000 0 0 $X=9232000 $Y=7056000
X4802 24 4692 ICV_9 $T=9296000 8912000 0 0 $X=9296000 $Y=8912000
X4803 24 4693 ICV_9 $T=9544000 1488000 0 0 $X=9544000 $Y=1488000
X4804 24 4694 ICV_9 $T=9544000 2880000 0 0 $X=9544000 $Y=2880000
X4805 24 4695 ICV_9 $T=9568000 96000 0 0 $X=9568000 $Y=96000
X4806 24 4696 ICV_9 $T=9600000 2416000 0 0 $X=9600000 $Y=2416000
X4807 24 4697 ICV_9 $T=9624000 3808000 0 0 $X=9624000 $Y=3808000
X4808 24 4698 ICV_9 $T=9632000 1952000 0 0 $X=9632000 $Y=1952000
X4809 24 4699 ICV_9 $T=9872000 96000 0 0 $X=9872000 $Y=96000
X4810 24 4700 ICV_9 $T=9880000 2880000 0 0 $X=9880000 $Y=2880000
X4811 24 4701 ICV_9 $T=9888000 9840000 0 0 $X=9888000 $Y=9840000
X4812 24 4702 ICV_9 $T=10008000 6128000 0 0 $X=10008000 $Y=6128000
X4813 24 4703 ICV_9 $T=10024000 12392000 0 0 $X=10024000 $Y=12392000
X4814 24 2351 ICV_9 $T=10080000 8216000 0 0 $X=10080000 $Y=8216000
X4815 24 4704 ICV_9 $T=10096000 1488000 0 0 $X=10096000 $Y=1488000
X4816 24 4705 ICV_9 $T=10136000 6592000 0 0 $X=10136000 $Y=6592000
X4817 24 4706 ICV_9 $T=10184000 9840000 0 0 $X=10184000 $Y=9840000
X4818 24 4707 ICV_9 $T=10216000 9376000 0 0 $X=10216000 $Y=9376000
X4819 24 4708 ICV_9 $T=10248000 7056000 0 0 $X=10248000 $Y=7056000
X4820 24 4709 ICV_9 $T=10352000 4968000 0 0 $X=10352000 $Y=4968000
X4821 24 4710 ICV_9 $T=10552000 12856000 0 0 $X=10552000 $Y=12856000
X4822 24 4711 ICV_9 $T=10744000 6592000 0 0 $X=10744000 $Y=6592000
X4823 24 4712 ICV_9 $T=10752000 7288000 0 0 $X=10752000 $Y=7288000
X4824 24 4713 ICV_9 $T=10784000 8680000 0 0 $X=10784000 $Y=8680000
X4825 24 4714 ICV_9 $T=10808000 4040000 0 0 $X=10808000 $Y=4040000
X4826 24 4715 ICV_9 $T=10880000 5432000 0 0 $X=10880000 $Y=5432000
X4827 24 4716 ICV_9 $T=10920000 10304000 0 0 $X=10920000 $Y=10304000
X4828 24 4717 ICV_9 $T=10976000 7056000 0 0 $X=10976000 $Y=7056000
X4829 24 4718 ICV_9 $T=11008000 8912000 0 0 $X=11008000 $Y=8912000
X4830 24 4719 ICV_9 $T=11008000 11000000 0 0 $X=11008000 $Y=11000000
X4831 24 4720 ICV_9 $T=11184000 5200000 0 0 $X=11184000 $Y=5200000
X4832 24 4103 ICV_9 $T=11256000 3344000 0 0 $X=11256000 $Y=3344000
X4833 24 4721 ICV_9 $T=11304000 7288000 0 0 $X=11304000 $Y=7288000
X4834 24 4722 ICV_9 $T=11312000 8912000 0 0 $X=11312000 $Y=8912000
X4835 24 4723 ICV_9 $T=11368000 6360000 0 0 $X=11368000 $Y=6360000
X4836 24 4724 ICV_9 $T=11488000 4040000 0 0 $X=11488000 $Y=4040000
X4837 24 4725 ICV_9 $T=11552000 7520000 0 0 $X=11552000 $Y=7520000
X4838 24 4726 ICV_9 $T=11720000 11232000 0 0 $X=11720000 $Y=11232000
X4839 24 4727 ICV_9 $T=11760000 11696000 0 0 $X=11760000 $Y=11696000
X4840 24 4728 ICV_9 $T=11800000 11464000 0 0 $X=11800000 $Y=11464000
X4841 24 4729 ICV_9 $T=11920000 4272000 0 0 $X=11920000 $Y=4272000
X4842 24 4730 ICV_9 $T=11928000 3344000 0 0 $X=11928000 $Y=3344000
X4843 24 4731 ICV_9 $T=11984000 4736000 0 0 $X=11984000 $Y=4736000
X4844 24 4732 ICV_9 $T=12040000 4968000 0 0 $X=12040000 $Y=4968000
X4845 24 4733 dff $T=152000 96000 0 0 $X=152000 $Y=96000
X4846 24 4734 dff $T=152000 328000 0 0 $X=152000 $Y=328000
X4847 24 4735 dff $T=152000 560000 0 0 $X=152000 $Y=560000
X4848 24 4736 dff $T=152000 792000 0 0 $X=152000 $Y=792000
X4849 24 4737 dff $T=152000 1024000 0 0 $X=152000 $Y=1024000
X4850 24 4738 dff $T=152000 1256000 0 0 $X=152000 $Y=1256000
X4851 24 4739 dff $T=152000 1488000 0 0 $X=152000 $Y=1488000
X4852 24 4740 dff $T=152000 1952000 0 0 $X=152000 $Y=1952000
X4853 24 4741 dff $T=152000 2184000 0 0 $X=152000 $Y=2184000
X4854 24 4742 dff $T=152000 2416000 0 0 $X=152000 $Y=2416000
X4855 24 4743 dff $T=152000 2880000 0 0 $X=152000 $Y=2880000
X4856 24 4744 dff $T=152000 4272000 0 0 $X=152000 $Y=4272000
X4857 24 4745 dff $T=184000 1720000 0 0 $X=184000 $Y=1720000
X4858 24 4746 dff $T=216000 3344000 0 0 $X=216000 $Y=3344000
X4859 24 4747 dff $T=376000 2648000 0 0 $X=376000 $Y=2648000
X4860 24 4748 dff $T=424000 2416000 0 0 $X=424000 $Y=2416000
X4861 24 4749 dff $T=440000 1952000 0 0 $X=440000 $Y=1952000
X4862 24 4750 dff $T=512000 328000 0 0 $X=512000 $Y=328000
X4863 24 4751 dff $T=560000 1256000 0 0 $X=560000 $Y=1256000
X4864 24 4752 dff $T=568000 792000 0 0 $X=568000 $Y=792000
X4865 24 4753 dff $T=568000 1488000 0 0 $X=568000 $Y=1488000
X4866 24 4754 dff $T=584000 1720000 0 0 $X=584000 $Y=1720000
X4867 24 4755 dff $T=782000 560000 1 180 $X=624000 $Y=560000
X4868 24 4756 dff $T=632000 2880000 0 0 $X=632000 $Y=2880000
X4869 24 4757 dff $T=822000 2648000 1 180 $X=664000 $Y=2648000
X4870 24 4758 dff $T=736000 3344000 0 0 $X=736000 $Y=3344000
X4871 24 4759 dff $T=966000 1720000 1 180 $X=808000 $Y=1720000
X4872 24 4760 dff $T=808000 2184000 0 0 $X=808000 $Y=2184000
X4873 24 4761 dff $T=856000 96000 0 0 $X=856000 $Y=96000
X4874 24 4762 dff $T=912000 1024000 0 0 $X=912000 $Y=1024000
X4875 24 4763 dff $T=1078000 328000 1 180 $X=920000 $Y=328000
X4876 24 4764 dff $T=928000 3344000 0 0 $X=928000 $Y=3344000
X4877 24 4765 dff $T=968000 2184000 0 0 $X=968000 $Y=2184000
X4878 24 4766 dff $T=976000 1256000 0 0 $X=976000 $Y=1256000
X4879 24 4767 dff $T=1150000 3576000 1 180 $X=992000 $Y=3576000
X4880 24 4768 dff $T=1190000 1952000 1 180 $X=1032000 $Y=1952000
X4881 24 4769 dff $T=1190000 3808000 1 180 $X=1032000 $Y=3808000
X4882 24 4770 dff $T=1040000 792000 0 0 $X=1040000 $Y=792000
X4883 24 4771 dff $T=1104000 2416000 0 0 $X=1104000 $Y=2416000
X4884 24 4772 dff $T=1112000 1488000 0 0 $X=1112000 $Y=1488000
X4885 24 4773 dff $T=1200000 1024000 0 0 $X=1200000 $Y=1024000
X4886 24 4774 dff $T=1208000 328000 0 0 $X=1208000 $Y=328000
X4887 24 4775 dff $T=1414000 96000 1 180 $X=1256000 $Y=96000
X4888 24 4776 dff $T=1430000 1488000 1 180 $X=1272000 $Y=1488000
X4889 24 4777 dff $T=1486000 560000 1 180 $X=1328000 $Y=560000
X4890 24 4778 dff $T=1486000 2416000 1 180 $X=1328000 $Y=2416000
X4891 24 4779 dff $T=1526000 328000 1 180 $X=1368000 $Y=328000
X4892 24 4780 dff $T=1384000 1720000 0 0 $X=1384000 $Y=1720000
X4893 24 4781 dff $T=1392000 1024000 0 0 $X=1392000 $Y=1024000
X4894 24 4782 dff $T=1566000 1952000 1 180 $X=1408000 $Y=1952000
X4895 24 4783 dff $T=1408000 3576000 0 0 $X=1408000 $Y=3576000
X4896 24 4784 dff $T=1536000 792000 0 0 $X=1536000 $Y=792000
X4897 24 4785 dff $T=1560000 2184000 0 0 $X=1560000 $Y=2184000
X4898 24 4786 dff $T=1766000 96000 1 180 $X=1608000 $Y=96000
X4899 24 4787 dff $T=1624000 2648000 0 0 $X=1624000 $Y=2648000
X4900 24 4788 dff $T=1648000 560000 0 0 $X=1648000 $Y=560000
X4901 24 4789 dff $T=1672000 1256000 0 0 $X=1672000 $Y=1256000
X4902 24 4790 dff $T=1680000 1024000 0 0 $X=1680000 $Y=1024000
X4903 24 4791 dff $T=1712000 1720000 0 0 $X=1712000 $Y=1720000
X4904 24 4792 dff $T=1720000 328000 0 0 $X=1720000 $Y=328000
X4905 24 4793 dff $T=1728000 2416000 0 0 $X=1728000 $Y=2416000
X4906 24 4794 dff $T=1950000 2184000 1 180 $X=1792000 $Y=2184000
X4907 24 4795 dff $T=1958000 3112000 1 180 $X=1800000 $Y=3112000
X4908 24 4796 dff $T=1990000 96000 1 180 $X=1832000 $Y=96000
X4909 24 4797 dff $T=1872000 560000 0 0 $X=1872000 $Y=560000
X4910 24 4798 dff $T=1872000 1720000 0 0 $X=1872000 $Y=1720000
X4911 24 4799 dff $T=1920000 1952000 0 0 $X=1920000 $Y=1952000
X4912 24 4800 dff $T=2102000 792000 1 180 $X=1944000 $Y=792000
X4913 24 4801 dff $T=1968000 1488000 0 0 $X=1968000 $Y=1488000
X4914 24 4802 dff $T=2016000 2880000 0 0 $X=2016000 $Y=2880000
X4915 24 4803 dff $T=2182000 2648000 1 180 $X=2024000 $Y=2648000
X4916 24 4804 dff $T=2104000 1024000 0 0 $X=2104000 $Y=1024000
X4917 24 4805 dff $T=2120000 96000 0 0 $X=2120000 $Y=96000
X4918 24 4806 dff $T=2286000 328000 1 180 $X=2128000 $Y=328000
X4919 24 4807 dff $T=2128000 2416000 0 0 $X=2128000 $Y=2416000
X4920 24 4808 dff $T=2144000 2184000 0 0 $X=2144000 $Y=2184000
X4921 24 4809 dff $T=2334000 2880000 1 180 $X=2176000 $Y=2880000
X4922 24 4810 dff $T=2350000 1720000 1 180 $X=2192000 $Y=1720000
X4923 24 4811 dff $T=2264000 6824000 0 0 $X=2264000 $Y=6824000
X4924 24 4812 dff $T=2272000 1256000 0 0 $X=2272000 $Y=1256000
X4925 24 4813 dff $T=2438000 1488000 1 180 $X=2280000 $Y=1488000
X4926 24 4814 dff $T=2296000 2648000 0 0 $X=2296000 $Y=2648000
X4927 24 4815 dff $T=2352000 792000 0 0 $X=2352000 $Y=792000
X4928 24 4816 dff $T=2400000 560000 0 0 $X=2400000 $Y=560000
X4929 24 4817 dff $T=2496000 2416000 0 0 $X=2496000 $Y=2416000
X4930 24 4818 dff $T=2670000 792000 1 180 $X=2512000 $Y=792000
X4931 24 4819 dff $T=2560000 1256000 0 0 $X=2560000 $Y=1256000
X4932 24 4820 dff $T=2734000 1024000 1 180 $X=2576000 $Y=1024000
X4933 24 4821 dff $T=2608000 1720000 0 0 $X=2608000 $Y=1720000
X4934 24 4822 dff $T=2616000 2648000 0 0 $X=2616000 $Y=2648000
X4935 24 4823 dff $T=2664000 328000 0 0 $X=2664000 $Y=328000
X4936 24 4824 dff $T=2744000 2880000 0 0 $X=2744000 $Y=2880000
X4937 24 4825 dff $T=2800000 792000 0 0 $X=2800000 $Y=792000
X4938 24 4826 dff $T=2816000 1952000 0 0 $X=2816000 $Y=1952000
X4939 24 4827 dff $T=2816000 6824000 0 0 $X=2816000 $Y=6824000
X4940 24 4828 dff $T=2864000 1024000 0 0 $X=2864000 $Y=1024000
X4941 24 4829 dff $T=3078000 2416000 1 180 $X=2920000 $Y=2416000
X4942 24 4830 dff $T=2936000 2648000 0 0 $X=2936000 $Y=2648000
X4943 24 4831 dff $T=2960000 2880000 0 0 $X=2960000 $Y=2880000
X4944 24 4832 dff $T=3198000 2184000 1 180 $X=3040000 $Y=2184000
X4945 24 4833 dff $T=3256000 96000 0 0 $X=3256000 $Y=96000
X4946 24 4834 dff $T=3264000 328000 0 0 $X=3264000 $Y=328000
X4947 24 4835 dff $T=3920000 96000 0 0 $X=3920000 $Y=96000
X4948 24 4836 dff $T=4494000 328000 1 180 $X=4336000 $Y=328000
X4949 24 4837 dff $T=4360000 96000 0 0 $X=4360000 $Y=96000
X4950 24 4838 dff $T=4718000 1488000 1 180 $X=4560000 $Y=1488000
X4951 24 2326 dff $T=6208000 96000 0 0 $X=6208000 $Y=96000
X4952 24 4839 dff $T=10542000 1488000 1 180 $X=10384000 $Y=1488000
X4953 24 4840 dff $T=10582000 1024000 1 180 $X=10424000 $Y=1024000
X4954 24 4841 dff $T=10568000 1256000 0 0 $X=10568000 $Y=1256000
X4955 24 4842 dff $T=10856000 1256000 0 0 $X=10856000 $Y=1256000
X4956 24 4843 dff $T=11046000 1488000 1 180 $X=10888000 $Y=1488000
X4957 24 4844 dff $T=11000000 560000 0 0 $X=11000000 $Y=560000
X4958 24 4845 dff $T=11286000 6824000 1 180 $X=11128000 $Y=6824000
X4959 24 4846 dff $T=11494000 6824000 1 180 $X=11336000 $Y=6824000
X4960 24 2357 dff $T=11520000 8680000 0 0 $X=11520000 $Y=8680000
X4961 24 4847 dff $T=11632000 1024000 0 0 $X=11632000 $Y=1024000
X4962 24 4848 dff $T=11648000 1720000 0 0 $X=11648000 $Y=1720000
X4963 24 4849 dff $T=11936000 6824000 0 0 $X=11936000 $Y=6824000
X4964 24 ICV_10 $T=1616000 8216000 0 0 $X=1616000 $Y=8216000
X4965 24 ICV_10 $T=1752000 6128000 0 0 $X=1752000 $Y=6128000
X4966 24 ICV_10 $T=2248000 3808000 0 0 $X=2248000 $Y=3808000
X4967 24 ICV_10 $T=2800000 3576000 0 0 $X=2800000 $Y=3576000
X4968 24 ICV_10 $T=3592000 9144000 0 0 $X=3592000 $Y=9144000
X4969 24 ICV_10 $T=3792000 2880000 0 0 $X=3792000 $Y=2880000
X4970 24 ICV_10 $T=4168000 6360000 0 0 $X=4168000 $Y=6360000
X4971 24 ICV_10 $T=4368000 2184000 0 0 $X=4368000 $Y=2184000
X4972 24 ICV_10 $T=4800000 11232000 0 0 $X=4800000 $Y=11232000
X4973 24 ICV_10 $T=5072000 2648000 0 0 $X=5072000 $Y=2648000
X4974 24 ICV_10 $T=5192000 6592000 0 0 $X=5192000 $Y=6592000
X4975 24 ICV_10 $T=5376000 2184000 0 0 $X=5376000 $Y=2184000
X4976 24 ICV_10 $T=5488000 12624000 0 0 $X=5488000 $Y=12624000
X4977 24 ICV_10 $T=5560000 560000 0 0 $X=5560000 $Y=560000
X4978 24 ICV_10 $T=6040000 3576000 0 0 $X=6040000 $Y=3576000
X4979 24 ICV_10 $T=6680000 7984000 0 0 $X=6680000 $Y=7984000
X4980 24 ICV_10 $T=6944000 12856000 0 0 $X=6944000 $Y=12856000
X4981 24 ICV_10 $T=7080000 1720000 0 0 $X=7080000 $Y=1720000
X4982 24 ICV_10 $T=7136000 4040000 0 0 $X=7136000 $Y=4040000
X4983 24 ICV_10 $T=7176000 8216000 0 0 $X=7176000 $Y=8216000
X4984 24 ICV_10 $T=8080000 6128000 0 0 $X=8080000 $Y=6128000
X4985 24 ICV_10 $T=8448000 8680000 0 0 $X=8448000 $Y=8680000
X4986 24 ICV_10 $T=9512000 328000 0 0 $X=9512000 $Y=328000
X4987 24 ICV_10 $T=9520000 2648000 0 0 $X=9520000 $Y=2648000
X4988 24 ICV_10 $T=10208000 10768000 0 0 $X=10208000 $Y=10768000
X4989 24 ICV_10 $T=10232000 8912000 0 0 $X=10232000 $Y=8912000
X4990 24 ICV_10 $T=10480000 4504000 0 0 $X=10480000 $Y=4504000
X4991 24 ICV_10 $T=10512000 10768000 0 0 $X=10512000 $Y=10768000
X4992 24 ICV_10 $T=10848000 10536000 0 0 $X=10848000 $Y=10536000
X4993 24 ICV_10 $T=11240000 5432000 0 0 $X=11240000 $Y=5432000
X4994 24 ICV_10 $T=11328000 3808000 0 0 $X=11328000 $Y=3808000
X4995 24 ICV_10 $T=11864000 3576000 0 0 $X=11864000 $Y=3576000
X4996 24 4850 and03 $T=232000 10072000 0 0 $X=232000 $Y=10072000
X4997 24 4851 and03 $T=305500 11928000 1 180 $X=256000 $Y=11928000
X4998 24 4852 and03 $T=337500 10072000 1 180 $X=288000 $Y=10072000
X4999 24 4853 and03 $T=361500 11928000 1 180 $X=312000 $Y=11928000
X5000 24 4854 and03 $T=344000 10072000 0 0 $X=344000 $Y=10072000
X5001 24 4855 and03 $T=368000 11928000 0 0 $X=368000 $Y=11928000
X5002 24 4856 and03 $T=449500 10072000 1 180 $X=400000 $Y=10072000
X5003 24 4857 and03 $T=456000 10072000 0 0 $X=456000 $Y=10072000
X5004 24 4858 and03 $T=521500 12392000 1 180 $X=472000 $Y=12392000
X5005 24 4859 and03 $T=504000 10768000 0 0 $X=504000 $Y=10768000
X5006 24 4860 and03 $T=577500 12392000 1 180 $X=528000 $Y=12392000
X5007 24 4861 and03 $T=633500 12392000 1 180 $X=584000 $Y=12392000
X5008 24 4862 and03 $T=616000 10072000 0 0 $X=616000 $Y=10072000
X5009 24 4863 and03 $T=729500 12160000 1 180 $X=680000 $Y=12160000
X5010 24 4864 and03 $T=753500 10768000 1 180 $X=704000 $Y=10768000
X5011 24 4865 and03 $T=753500 11000000 1 180 $X=704000 $Y=11000000
X5012 24 4866 and03 $T=753500 11232000 1 180 $X=704000 $Y=11232000
X5013 24 4867 and03 $T=785500 12160000 1 180 $X=736000 $Y=12160000
X5014 24 4868 and03 $T=809500 10768000 1 180 $X=760000 $Y=10768000
X5015 24 4869 and03 $T=809500 11232000 1 180 $X=760000 $Y=11232000
X5016 24 4870 and03 $T=768000 11464000 0 0 $X=768000 $Y=11464000
X5017 24 4871 and03 $T=841500 11000000 1 180 $X=792000 $Y=11000000
X5018 24 4872 and03 $T=865500 10768000 1 180 $X=816000 $Y=10768000
X5019 24 4873 and03 $T=848000 11000000 0 0 $X=848000 $Y=11000000
X5020 24 4874 and03 $T=905500 10304000 1 180 $X=856000 $Y=10304000
X5021 24 4875 and03 $T=872000 10768000 0 0 $X=872000 $Y=10768000
X5022 24 4876 and03 $T=872000 11232000 0 0 $X=872000 $Y=11232000
X5023 24 4877 and03 $T=937500 12392000 1 180 $X=888000 $Y=12392000
X5024 24 4878 and03 $T=904000 10072000 0 0 $X=904000 $Y=10072000
X5025 24 4879 and03 $T=961500 10304000 1 180 $X=912000 $Y=10304000
X5026 24 4880 and03 $T=977500 10768000 1 180 $X=928000 $Y=10768000
X5027 24 4881 and03 $T=944000 12160000 0 0 $X=944000 $Y=12160000
X5028 24 4882 and03 $T=1000000 10072000 0 0 $X=1000000 $Y=10072000
X5029 24 4883 and03 $T=1057500 12392000 1 180 $X=1008000 $Y=12392000
X5030 24 4884 and03 $T=1073500 10768000 1 180 $X=1024000 $Y=10768000
X5031 24 4885 and03 $T=1113500 12392000 1 180 $X=1064000 $Y=12392000
X5032 24 4886 and03 $T=1129500 10768000 1 180 $X=1080000 $Y=10768000
X5033 24 4887 and03 $T=1161500 11928000 1 180 $X=1112000 $Y=11928000
X5034 24 4888 and03 $T=1169500 12392000 1 180 $X=1120000 $Y=12392000
X5035 24 4889 and03 $T=1185500 10768000 1 180 $X=1136000 $Y=10768000
X5036 24 4890 and03 $T=1201500 11000000 1 180 $X=1152000 $Y=11000000
X5037 24 4891 and03 $T=1209500 10536000 1 180 $X=1160000 $Y=10536000
X5038 24 4892 and03 $T=1200000 10072000 0 0 $X=1200000 $Y=10072000
X5039 24 4893 and03 $T=1257500 11000000 1 180 $X=1208000 $Y=11000000
X5040 24 2299 and03 $T=1265500 10304000 1 180 $X=1216000 $Y=10304000
X5041 24 4894 and03 $T=1224000 10768000 0 0 $X=1224000 $Y=10768000
X5042 24 4895 and03 $T=1272000 10304000 0 0 $X=1272000 $Y=10304000
X5043 24 4896 and03 $T=1280000 10768000 0 0 $X=1280000 $Y=10768000
X5044 24 4897 and03 $T=1336000 10768000 0 0 $X=1336000 $Y=10768000
X5045 24 4898 and03 $T=1392000 10768000 0 0 $X=1392000 $Y=10768000
X5046 24 4899 and03 $T=1448000 10768000 0 0 $X=1448000 $Y=10768000
X5047 24 4900 and03 $T=1553500 10768000 1 180 $X=1504000 $Y=10768000
X5048 24 4901 and03 $T=1553500 11928000 1 180 $X=1504000 $Y=11928000
X5049 24 4902 and03 $T=1609500 10768000 1 180 $X=1560000 $Y=10768000
X5050 24 4903 and03 $T=1609500 11928000 1 180 $X=1560000 $Y=11928000
X5051 24 4904 and03 $T=1592000 10536000 0 0 $X=1592000 $Y=10536000
X5052 24 4905 and03 $T=2048000 10304000 0 0 $X=2048000 $Y=10304000
X5053 24 4906 and03 $T=2208000 10304000 0 0 $X=2208000 $Y=10304000
X5054 24 4907 and03 $T=2264000 10304000 0 0 $X=2264000 $Y=10304000
X5055 24 4908 and03 $T=2360000 10304000 0 0 $X=2360000 $Y=10304000
X5056 24 4909 and03 $T=2456000 10304000 0 0 $X=2456000 $Y=10304000
X5057 24 4910 and03 $T=2512000 10304000 0 0 $X=2512000 $Y=10304000
X5058 24 4911 and03 $T=2568000 10304000 0 0 $X=2568000 $Y=10304000
X5059 24 4912 and03 $T=3016000 10304000 0 0 $X=3016000 $Y=10304000
X5060 24 4913 and03 $T=3072000 10304000 0 0 $X=3072000 $Y=10304000
X5061 24 4914 and03 $T=3456000 10072000 0 0 $X=3456000 $Y=10072000
X5062 24 4915 and03 $T=3552000 10072000 0 0 $X=3552000 $Y=10072000
X5063 24 4916 and03 $T=3608000 10072000 0 0 $X=3608000 $Y=10072000
X5064 24 4917 and03 $T=3760000 10304000 0 0 $X=3760000 $Y=10304000
X5065 24 4918 and03 $T=3848000 10304000 0 0 $X=3848000 $Y=10304000
X5066 24 4919 and03 $T=3944000 10304000 0 0 $X=3944000 $Y=10304000
X5067 24 4920 and03 $T=4000000 10304000 0 0 $X=4000000 $Y=10304000
X5068 24 4921 and03 $T=4393500 10304000 1 180 $X=4344000 $Y=10304000
X5069 24 4922 and03 $T=4400000 10304000 0 0 $X=4400000 $Y=10304000
X5070 24 4923 and03 $T=4456000 10304000 0 0 $X=4456000 $Y=10304000
X5071 24 4924 and03 $T=4512000 10304000 0 0 $X=4512000 $Y=10304000
X5072 24 4925 and03 $T=4617500 10304000 1 180 $X=4568000 $Y=10304000
X5073 24 4926 and03 $T=4681500 10536000 1 180 $X=4632000 $Y=10536000
X5074 24 4927 and03 $T=4664000 10304000 0 0 $X=4664000 $Y=10304000
X5075 24 4928 and03 $T=4688000 10536000 0 0 $X=4688000 $Y=10536000
X5076 24 4929 and03 $T=4744000 10536000 0 0 $X=4744000 $Y=10536000
X5077 24 4930 and03 $T=5040000 10304000 0 0 $X=5040000 $Y=10304000
X5078 24 4931 and03 $T=5072000 10768000 0 0 $X=5072000 $Y=10768000
X5079 24 4932 and03 $T=5177500 10304000 1 180 $X=5128000 $Y=10304000
X5080 24 4933 and03 $T=5128000 10768000 0 0 $X=5128000 $Y=10768000
X5081 24 4934 and03 $T=5152000 10536000 0 0 $X=5152000 $Y=10536000
X5082 24 4935 and03 $T=5152000 11000000 0 0 $X=5152000 $Y=11000000
X5083 24 4936 and03 $T=5184000 10304000 0 0 $X=5184000 $Y=10304000
X5084 24 4937 and03 $T=5184000 10768000 0 0 $X=5184000 $Y=10768000
X5085 24 4938 and03 $T=5232000 11232000 0 0 $X=5232000 $Y=11232000
X5086 24 4939 and03 $T=5240000 10768000 0 0 $X=5240000 $Y=10768000
X5087 24 4940 and03 $T=5248000 10536000 0 0 $X=5248000 $Y=10536000
X5088 24 4941 and03 $T=5280000 10304000 0 0 $X=5280000 $Y=10304000
X5089 24 4942 and03 $T=5312000 11000000 0 0 $X=5312000 $Y=11000000
X5090 24 4943 and03 $T=5336000 10304000 0 0 $X=5336000 $Y=10304000
X5091 24 4944 and03 $T=5504000 10304000 0 0 $X=5504000 $Y=10304000
X5092 24 4945 and03 $T=5648000 10536000 0 0 $X=5648000 $Y=10536000
X5093 24 4946 and03 $T=5793500 11000000 1 180 $X=5744000 $Y=11000000
X5094 24 4947 and03 $T=5752000 11232000 0 0 $X=5752000 $Y=11232000
X5095 24 4948 and03 $T=5832000 11000000 0 0 $X=5832000 $Y=11000000
X5096 24 4949 and03 $T=5880000 10304000 0 0 $X=5880000 $Y=10304000
X5097 24 4950 and03 $T=5880000 11464000 0 0 $X=5880000 $Y=11464000
X5098 24 4951 and03 $T=5888000 11000000 0 0 $X=5888000 $Y=11000000
X5099 24 4952 and03 $T=5912000 11232000 0 0 $X=5912000 $Y=11232000
X5100 24 4953 and03 $T=5936000 10304000 0 0 $X=5936000 $Y=10304000
X5101 24 4954 and03 $T=5944000 11000000 0 0 $X=5944000 $Y=11000000
X5102 24 4955 and03 $T=5992000 10304000 0 0 $X=5992000 $Y=10304000
X5103 24 4956 and03 $T=6048000 10304000 0 0 $X=6048000 $Y=10304000
X5104 24 4957 and03 $T=7304000 11928000 0 0 $X=7304000 $Y=11928000
X5105 24 4958 and03 $T=7409500 11928000 1 180 $X=7360000 $Y=11928000
X5106 24 4959 and03 $T=7497500 11928000 1 180 $X=7448000 $Y=11928000
X5107 24 4960 and03 $T=7873500 11928000 1 180 $X=7824000 $Y=11928000
X5108 24 4961 and03 $T=7848000 11696000 0 0 $X=7848000 $Y=11696000
X5109 24 4962 and03 $T=7904000 11696000 0 0 $X=7904000 $Y=11696000
X5110 24 4963 and03 $T=8937500 11696000 1 180 $X=8888000 $Y=11696000
X5111 24 4964 and03 $T=8961500 11928000 1 180 $X=8912000 $Y=11928000
X5112 24 4100 and03 $T=8920000 11464000 0 0 $X=8920000 $Y=11464000
X5113 24 4965 and03 $T=9016000 11928000 0 0 $X=9016000 $Y=11928000
X5114 24 4966 and03 $T=9136000 11232000 0 0 $X=9136000 $Y=11232000
X5115 24 4967 and03 $T=9176000 11464000 0 0 $X=9176000 $Y=11464000
X5116 24 4968 and03 $T=9353500 11464000 1 180 $X=9304000 $Y=11464000
X5117 24 4969 and03 $T=9409500 11464000 1 180 $X=9360000 $Y=11464000
X5118 24 4970 and03 $T=9473500 12624000 1 180 $X=9424000 $Y=12624000
X5119 24 4971 and03 $T=9489500 12856000 1 180 $X=9440000 $Y=12856000
X5120 24 4972 and03 $T=9480000 12624000 0 0 $X=9480000 $Y=12624000
X5121 24 4973 and03 $T=9528000 13088000 0 0 $X=9528000 $Y=13088000
X5122 24 4974 and03 $T=9585500 12624000 1 180 $X=9536000 $Y=12624000
X5123 24 4975 and03 $T=9576000 12856000 0 0 $X=9576000 $Y=12856000
X5124 24 4976 and03 $T=9592000 12624000 0 0 $X=9592000 $Y=12624000
X5125 24 4977 and03 $T=9673500 13088000 1 180 $X=9624000 $Y=13088000
X5126 24 4978 and03 $T=9681500 12856000 1 180 $X=9632000 $Y=12856000
X5127 24 4979 and03 $T=9648000 12624000 0 0 $X=9648000 $Y=12624000
X5128 24 4980 and03 $T=9704000 12624000 0 0 $X=9704000 $Y=12624000
X5129 24 4981 and03 $T=9785500 11928000 1 180 $X=9736000 $Y=11928000
X5130 24 4982 and03 $T=9760000 12624000 0 0 $X=9760000 $Y=12624000
X5131 24 4983 and03 $T=9760000 13088000 0 0 $X=9760000 $Y=13088000
X5132 24 4984 and03 $T=9817500 12856000 1 180 $X=9768000 $Y=12856000
X5133 24 4985 and03 $T=9792000 11928000 0 0 $X=9792000 $Y=11928000
X5134 24 4986 and03 $T=9865500 13088000 1 180 $X=9816000 $Y=13088000
X5135 24 4987 and03 $T=9873500 12856000 1 180 $X=9824000 $Y=12856000
X5136 24 4988 and03 $T=9832000 11464000 0 0 $X=9832000 $Y=11464000
X5137 24 4989 and03 $T=9921500 13088000 1 180 $X=9872000 $Y=13088000
X5138 24 4990 and03 $T=9945500 11696000 1 180 $X=9896000 $Y=11696000
X5139 24 4991 and03 $T=9896000 12624000 0 0 $X=9896000 $Y=12624000
X5140 24 4992 and03 $T=9912000 12856000 0 0 $X=9912000 $Y=12856000
X5141 24 4993 and03 $T=10025500 12160000 1 180 $X=9976000 $Y=12160000
X5142 24 4994 and03 $T=9984000 11696000 0 0 $X=9984000 $Y=11696000
X5143 24 4995 and03 $T=10049500 13088000 1 180 $X=10000000 $Y=13088000
X5144 24 4996 and03 $T=10024000 12624000 0 0 $X=10024000 $Y=12624000
X5145 24 4997 and03 $T=10040000 12856000 0 0 $X=10040000 $Y=12856000
X5146 24 4998 and03 $T=10056000 13088000 0 0 $X=10056000 $Y=13088000
X5147 24 4999 and03 $T=10145500 12856000 1 180 $X=10096000 $Y=12856000
X5148 24 5000 and03 $T=10112000 12624000 0 0 $X=10112000 $Y=12624000
X5149 24 5001 and03 $T=10112000 13088000 0 0 $X=10112000 $Y=13088000
X5150 24 5002 and03 $T=10152000 12856000 0 0 $X=10152000 $Y=12856000
X5151 24 5003 and03 $T=10168000 12624000 0 0 $X=10168000 $Y=12624000
X5152 24 5004 and03 $T=10273500 12624000 1 180 $X=10224000 $Y=12624000
X5153 24 5005 and03 $T=10289500 12856000 1 180 $X=10240000 $Y=12856000
X5154 24 5006 and03 $T=10289500 13088000 1 180 $X=10240000 $Y=13088000
X5155 24 5007 and03 $T=10280000 12624000 0 0 $X=10280000 $Y=12624000
X5156 24 5008 and03 $T=10336000 11696000 0 0 $X=10336000 $Y=11696000
X5157 24 5009 and03 $T=10745500 11696000 1 180 $X=10696000 $Y=11696000
X5158 24 5010 and03 $T=10777500 13088000 1 180 $X=10728000 $Y=13088000
X5159 24 5011 and03 $T=10752000 11696000 0 0 $X=10752000 $Y=11696000
X5160 24 5012 and03 $T=10848000 12856000 0 0 $X=10848000 $Y=12856000
X5161 24 5013 and03 $T=10945500 13088000 1 180 $X=10896000 $Y=13088000
X5162 24 5014 and03 $T=10953500 12856000 1 180 $X=10904000 $Y=12856000
X5163 24 5015 and03 $T=11009500 12856000 1 180 $X=10960000 $Y=12856000
X5164 24 5016 and03 $T=10992000 11696000 0 0 $X=10992000 $Y=11696000
X5165 24 5017 and03 $T=10992000 12160000 0 0 $X=10992000 $Y=12160000
X5166 24 5018 and03 $T=11048000 11696000 0 0 $X=11048000 $Y=11696000
X5167 24 5019 and03 $T=11080000 13320000 0 0 $X=11080000 $Y=13320000
X5168 24 5020 and03 $T=11104000 11696000 0 0 $X=11104000 $Y=11696000
X5169 24 5021 and03 $T=11168000 13320000 0 0 $X=11168000 $Y=13320000
X5170 24 5022 and03 $T=11184000 12624000 0 0 $X=11184000 $Y=12624000
X5171 24 5023 and03 $T=11200000 13552000 0 0 $X=11200000 $Y=13552000
X5172 24 5024 and03 $T=11224000 13320000 0 0 $X=11224000 $Y=13320000
X5173 24 5025 and03 $T=11312000 13320000 0 0 $X=11312000 $Y=13320000
X5174 24 5026 and03 $T=11544000 13088000 0 0 $X=11544000 $Y=13088000
X5175 24 5027 and03 $T=11592000 12856000 0 0 $X=11592000 $Y=12856000
X5176 24 5028 and03 $T=11728000 12160000 0 0 $X=11728000 $Y=12160000
X5177 24 5029 and03 $T=11792000 12160000 0 0 $X=11792000 $Y=12160000
X5178 24 5030 and03 $T=11800000 12856000 0 0 $X=11800000 $Y=12856000
X5179 24 5031 and03 $T=11848000 12160000 0 0 $X=11848000 $Y=12160000
X5180 24 5032 and03 $T=11856000 12856000 0 0 $X=11856000 $Y=12856000
X5181 24 5033 ICV_11 $T=1656000 5200000 0 0 $X=1656000 $Y=5200000
X5182 24 5034 ICV_11 $T=1672000 9840000 0 0 $X=1672000 $Y=9840000
X5183 24 5035 ICV_11 $T=1800000 6824000 0 0 $X=1800000 $Y=6824000
X5184 24 5036 ICV_11 $T=1928000 3344000 0 0 $X=1928000 $Y=3344000
X5185 24 5037 ICV_11 $T=1968000 5664000 0 0 $X=1968000 $Y=5664000
X5186 24 5038 ICV_11 $T=2352000 11000000 0 0 $X=2352000 $Y=11000000
X5187 24 5039 ICV_11 $T=2392000 13552000 0 0 $X=2392000 $Y=13552000
X5188 24 5040 ICV_11 $T=2656000 7752000 0 0 $X=2656000 $Y=7752000
X5189 24 5041 ICV_11 $T=2720000 8216000 0 0 $X=2720000 $Y=8216000
X5190 24 5042 ICV_11 $T=2936000 13552000 0 0 $X=2936000 $Y=13552000
X5191 24 5043 ICV_11 $T=2984000 12624000 0 0 $X=2984000 $Y=12624000
X5192 24 5044 ICV_11 $T=2992000 13088000 0 0 $X=2992000 $Y=13088000
X5193 24 5045 ICV_11 $T=3744000 2648000 0 0 $X=3744000 $Y=2648000
X5194 24 5046 ICV_11 $T=3808000 3112000 0 0 $X=3808000 $Y=3112000
X5195 24 5047 ICV_11 $T=3992000 5200000 0 0 $X=3992000 $Y=5200000
X5196 24 5048 ICV_11 $T=4232000 8216000 0 0 $X=4232000 $Y=8216000
X5197 24 5049 ICV_11 $T=4528000 13552000 0 0 $X=4528000 $Y=13552000
X5198 24 5050 ICV_11 $T=4776000 6824000 0 0 $X=4776000 $Y=6824000
X5199 24 5051 ICV_11 $T=4888000 5200000 0 0 $X=4888000 $Y=5200000
X5200 24 5052 ICV_11 $T=5080000 4504000 0 0 $X=5080000 $Y=4504000
X5201 24 5053 ICV_11 $T=5408000 3112000 0 0 $X=5408000 $Y=3112000
X5202 24 5054 ICV_11 $T=5440000 8912000 0 0 $X=5440000 $Y=8912000
X5203 24 5055 ICV_11 $T=5488000 1024000 0 0 $X=5488000 $Y=1024000
X5204 24 5056 ICV_11 $T=5520000 4272000 0 0 $X=5520000 $Y=4272000
X5205 24 5057 ICV_11 $T=5528000 3344000 0 0 $X=5528000 $Y=3344000
X5206 24 5058 ICV_11 $T=5600000 10072000 0 0 $X=5600000 $Y=10072000
X5207 24 5059 ICV_11 $T=5800000 5432000 0 0 $X=5800000 $Y=5432000
X5208 24 5060 ICV_11 $T=5824000 13552000 0 0 $X=5824000 $Y=13552000
X5209 24 5061 ICV_11 $T=5888000 6360000 0 0 $X=5888000 $Y=6360000
X5210 24 5062 ICV_11 $T=5968000 13088000 0 0 $X=5968000 $Y=13088000
X5211 24 5063 ICV_11 $T=6064000 8216000 0 0 $X=6064000 $Y=8216000
X5212 24 5064 ICV_11 $T=7256000 1488000 0 0 $X=7256000 $Y=1488000
X5213 24 5065 ICV_11 $T=7264000 4968000 0 0 $X=7264000 $Y=4968000
X5214 24 5066 ICV_11 $T=7304000 12856000 0 0 $X=7304000 $Y=12856000
X5215 24 5067 ICV_11 $T=7512000 11232000 0 0 $X=7512000 $Y=11232000
X5216 24 5068 ICV_11 $T=7528000 7288000 0 0 $X=7528000 $Y=7288000
X5217 24 5069 ICV_11 $T=7960000 12624000 0 0 $X=7960000 $Y=12624000
X5218 24 5070 ICV_11 $T=7968000 7056000 0 0 $X=7968000 $Y=7056000
X5219 24 5071 ICV_11 $T=9184000 8448000 0 0 $X=9184000 $Y=8448000
X5220 24 5072 ICV_11 $T=9256000 5432000 0 0 $X=9256000 $Y=5432000
X5221 24 5073 ICV_11 $T=9296000 11232000 0 0 $X=9296000 $Y=11232000
X5222 24 5074 ICV_11 $T=9408000 5200000 0 0 $X=9408000 $Y=5200000
X5223 24 5075 ICV_11 $T=9720000 560000 0 0 $X=9720000 $Y=560000
X5224 24 5076 ICV_11 $T=9800000 7752000 0 0 $X=9800000 $Y=7752000
X5225 24 5077 ICV_11 $T=9936000 4272000 0 0 $X=9936000 $Y=4272000
X5226 24 5078 ICV_11 $T=10008000 4736000 0 0 $X=10008000 $Y=4736000
X5227 24 5079 ICV_11 $T=10200000 7288000 0 0 $X=10200000 $Y=7288000
X5228 24 5080 ICV_11 $T=10200000 7520000 0 0 $X=10200000 $Y=7520000
X5229 24 5081 ICV_11 $T=10232000 6360000 0 0 $X=10232000 $Y=6360000
X5230 24 5082 ICV_11 $T=10392000 5664000 0 0 $X=10392000 $Y=5664000
X5231 24 5083 ICV_11 $T=10744000 2416000 0 0 $X=10744000 $Y=2416000
X5232 24 5084 ICV_11 $T=10808000 4272000 0 0 $X=10808000 $Y=4272000
X5233 24 5085 ICV_11 $T=10832000 9840000 0 0 $X=10832000 $Y=9840000
X5234 24 5086 ICV_11 $T=10920000 10768000 0 0 $X=10920000 $Y=10768000
X5235 24 5087 ICV_11 $T=11168000 11232000 0 0 $X=11168000 $Y=11232000
X5236 24 5088 ICV_11 $T=11288000 8448000 0 0 $X=11288000 $Y=8448000
X5237 24 5089 ICV_11 $T=11416000 8216000 0 0 $X=11416000 $Y=8216000
X5238 24 5090 ICV_11 $T=11560000 9840000 0 0 $X=11560000 $Y=9840000
X5239 24 5091 ICV_11 $T=11744000 8912000 0 0 $X=11744000 $Y=8912000
X5240 24 5092 ICV_11 $T=11784000 10768000 0 0 $X=11784000 $Y=10768000
X5241 24 5093 ICV_11 $T=11784000 11928000 0 0 $X=11784000 $Y=11928000
X5242 24 5094 ICV_11 $T=11792000 1952000 0 0 $X=11792000 $Y=1952000
X5243 24 5095 ICV_11 $T=11848000 5200000 0 0 $X=11848000 $Y=5200000
X5244 24 5096 ICV_11 $T=11848000 7752000 0 0 $X=11848000 $Y=7752000
X5245 24 ICV_12 $T=216000 10768000 0 0 $X=216000 $Y=10768000
X5246 24 ICV_12 $T=216000 12624000 0 0 $X=216000 $Y=12624000
X5247 24 ICV_12 $T=440000 11464000 0 0 $X=440000 $Y=11464000
X5248 24 ICV_12 $T=1344000 11696000 0 0 $X=1344000 $Y=11696000
X5249 24 ICV_12 $T=1888000 13552000 0 0 $X=1888000 $Y=13552000
X5250 24 ICV_12 $T=2792000 10304000 0 0 $X=2792000 $Y=10304000
X5251 24 ICV_12 $T=5400000 9840000 0 0 $X=5400000 $Y=9840000
X5252 24 ICV_12 $T=5616000 13320000 0 0 $X=5616000 $Y=13320000
X5253 24 ICV_12 $T=8312000 11928000 0 0 $X=8312000 $Y=11928000
X5254 24 ICV_12 $T=8688000 10072000 0 0 $X=8688000 $Y=10072000
X5255 24 ICV_12 $T=9584000 8680000 0 0 $X=9584000 $Y=8680000
X5256 24 ICV_12 $T=10176000 12160000 0 0 $X=10176000 $Y=12160000
X5257 24 ICV_12 $T=10488000 9840000 0 0 $X=10488000 $Y=9840000
X5258 24 ICV_12 $T=10944000 10072000 0 0 $X=10944000 $Y=10072000
X5259 24 ICV_12 $T=11832000 13552000 0 0 $X=11832000 $Y=13552000
X5260 24 5097 ICV_13 $T=1128000 11696000 0 0 $X=1128000 $Y=11696000
X5261 24 5098 ICV_13 $T=1648000 3344000 0 0 $X=1648000 $Y=3344000
X5262 24 5099 ICV_13 $T=1752000 7056000 0 0 $X=1752000 $Y=7056000
X5263 24 5100 ICV_13 $T=1768000 10304000 0 0 $X=1768000 $Y=10304000
X5264 24 5101 ICV_13 $T=1816000 10536000 0 0 $X=1816000 $Y=10536000
X5265 24 5102 ICV_13 $T=2024000 7520000 0 0 $X=2024000 $Y=7520000
X5266 24 5103 ICV_13 $T=2032000 9608000 0 0 $X=2032000 $Y=9608000
X5267 24 5104 ICV_13 $T=2272000 4272000 0 0 $X=2272000 $Y=4272000
X5268 24 5105 ICV_13 $T=2296000 8448000 0 0 $X=2296000 $Y=8448000
X5269 24 5106 ICV_13 $T=2776000 4040000 0 0 $X=2776000 $Y=4040000
X5270 24 5107 ICV_13 $T=3176000 5200000 0 0 $X=3176000 $Y=5200000
X5271 24 5108 ICV_13 $T=3192000 10304000 0 0 $X=3192000 $Y=10304000
X5272 24 5109 ICV_13 $T=3208000 4968000 0 0 $X=3208000 $Y=4968000
X5273 24 5110 ICV_13 $T=3264000 7288000 0 0 $X=3264000 $Y=7288000
X5274 24 5111 ICV_13 $T=3480000 12624000 0 0 $X=3480000 $Y=12624000
X5275 24 5112 ICV_13 $T=3632000 6824000 0 0 $X=3632000 $Y=6824000
X5276 24 5113 ICV_13 $T=3736000 10536000 0 0 $X=3736000 $Y=10536000
X5277 24 5114 ICV_13 $T=4088000 8448000 0 0 $X=4088000 $Y=8448000
X5278 24 5115 ICV_13 $T=4152000 10768000 0 0 $X=4152000 $Y=10768000
X5279 24 5116 ICV_13 $T=4472000 11696000 0 0 $X=4472000 $Y=11696000
X5280 24 5117 ICV_13 $T=4480000 11000000 0 0 $X=4480000 $Y=11000000
X5281 24 5118 ICV_13 $T=4544000 560000 0 0 $X=4544000 $Y=560000
X5282 24 5119 ICV_13 $T=4600000 12856000 0 0 $X=4600000 $Y=12856000
X5283 24 5120 ICV_13 $T=4944000 3808000 0 0 $X=4944000 $Y=3808000
X5284 24 5121 ICV_13 $T=5144000 9608000 0 0 $X=5144000 $Y=9608000
X5285 24 5122 ICV_13 $T=5160000 1720000 0 0 $X=5160000 $Y=1720000
X5286 24 5123 ICV_13 $T=5232000 1952000 0 0 $X=5232000 $Y=1952000
X5287 24 5124 ICV_13 $T=5440000 8680000 0 0 $X=5440000 $Y=8680000
X5288 24 5125 ICV_13 $T=5648000 13088000 0 0 $X=5648000 $Y=13088000
X5289 24 5126 ICV_13 $T=5720000 7984000 0 0 $X=5720000 $Y=7984000
X5290 24 5127 ICV_13 $T=5752000 8680000 0 0 $X=5752000 $Y=8680000
X5291 24 5128 ICV_13 $T=5768000 3808000 0 0 $X=5768000 $Y=3808000
X5292 24 5129 ICV_13 $T=5872000 12160000 0 0 $X=5872000 $Y=12160000
X5293 24 5130 ICV_13 $T=5936000 8448000 0 0 $X=5936000 $Y=8448000
X5294 24 5131 ICV_13 $T=6000000 3112000 0 0 $X=6000000 $Y=3112000
X5295 24 5132 ICV_13 $T=6048000 2648000 0 0 $X=6048000 $Y=2648000
X5296 24 5133 ICV_13 $T=6096000 2880000 0 0 $X=6096000 $Y=2880000
X5297 24 5134 ICV_13 $T=6184000 8912000 0 0 $X=6184000 $Y=8912000
X5298 24 5135 ICV_13 $T=6192000 12392000 0 0 $X=6192000 $Y=12392000
X5299 24 5136 ICV_13 $T=6272000 8680000 0 0 $X=6272000 $Y=8680000
X5300 24 5137 ICV_13 $T=6392000 12856000 0 0 $X=6392000 $Y=12856000
X5301 24 5138 ICV_13 $T=6704000 4736000 0 0 $X=6704000 $Y=4736000
X5302 24 5139 ICV_13 $T=6736000 4504000 0 0 $X=6736000 $Y=4504000
X5303 24 5140 ICV_13 $T=6744000 8680000 0 0 $X=6744000 $Y=8680000
X5304 24 5141 ICV_13 $T=6800000 4968000 0 0 $X=6800000 $Y=4968000
X5305 24 5142 ICV_13 $T=6800000 10072000 0 0 $X=6800000 $Y=10072000
X5306 24 5143 ICV_13 $T=6960000 6824000 0 0 $X=6960000 $Y=6824000
X5307 24 5144 ICV_13 $T=7040000 13320000 0 0 $X=7040000 $Y=13320000
X5308 24 5145 ICV_13 $T=7056000 3808000 0 0 $X=7056000 $Y=3808000
X5309 24 5146 ICV_13 $T=7080000 11000000 0 0 $X=7080000 $Y=11000000
X5310 24 5147 ICV_13 $T=7144000 8680000 0 0 $X=7144000 $Y=8680000
X5311 24 5148 ICV_13 $T=7256000 5432000 0 0 $X=7256000 $Y=5432000
X5312 24 5149 ICV_13 $T=7592000 560000 0 0 $X=7592000 $Y=560000
X5313 24 5150 ICV_13 $T=7592000 9608000 0 0 $X=7592000 $Y=9608000
X5314 24 5151 ICV_13 $T=7632000 10072000 0 0 $X=7632000 $Y=10072000
X5315 24 5152 ICV_13 $T=7704000 7984000 0 0 $X=7704000 $Y=7984000
X5316 24 5153 ICV_13 $T=7768000 6128000 0 0 $X=7768000 $Y=6128000
X5317 24 5154 ICV_13 $T=7800000 13320000 0 0 $X=7800000 $Y=13320000
X5318 24 5155 ICV_13 $T=7808000 5896000 0 0 $X=7808000 $Y=5896000
X5319 24 5156 ICV_13 $T=7848000 6360000 0 0 $X=7848000 $Y=6360000
X5320 24 5157 ICV_13 $T=7904000 4736000 0 0 $X=7904000 $Y=4736000
X5321 24 5158 ICV_13 $T=7936000 5200000 0 0 $X=7936000 $Y=5200000
X5322 24 5159 ICV_13 $T=8016000 560000 0 0 $X=8016000 $Y=560000
X5323 24 5160 ICV_13 $T=8176000 328000 0 0 $X=8176000 $Y=328000
X5324 24 5161 ICV_13 $T=8240000 4504000 0 0 $X=8240000 $Y=4504000
X5325 24 5162 ICV_13 $T=8320000 8448000 0 0 $X=8320000 $Y=8448000
X5326 24 5163 ICV_13 $T=8328000 5200000 0 0 $X=8328000 $Y=5200000
X5327 24 5164 ICV_13 $T=8352000 11232000 0 0 $X=8352000 $Y=11232000
X5328 24 5165 ICV_13 $T=8472000 1024000 0 0 $X=8472000 $Y=1024000
X5329 24 5166 ICV_13 $T=8528000 7752000 0 0 $X=8528000 $Y=7752000
X5330 24 5167 ICV_13 $T=8736000 1488000 0 0 $X=8736000 $Y=1488000
X5331 24 5168 ICV_13 $T=8744000 2648000 0 0 $X=8744000 $Y=2648000
X5332 24 5169 ICV_13 $T=8872000 7752000 0 0 $X=8872000 $Y=7752000
X5333 24 5170 ICV_13 $T=9016000 1488000 0 0 $X=9016000 $Y=1488000
X5334 24 5171 ICV_13 $T=9120000 9144000 0 0 $X=9120000 $Y=9144000
X5335 24 5172 ICV_13 $T=9232000 11928000 0 0 $X=9232000 $Y=11928000
X5336 24 5173 ICV_13 $T=9256000 10072000 0 0 $X=9256000 $Y=10072000
X5337 24 5174 ICV_13 $T=9416000 5664000 0 0 $X=9416000 $Y=5664000
X5338 24 5175 ICV_13 $T=9440000 3344000 0 0 $X=9440000 $Y=3344000
X5339 24 5176 ICV_13 $T=9536000 6592000 0 0 $X=9536000 $Y=6592000
X5340 24 5177 ICV_13 $T=9560000 2184000 0 0 $X=9560000 $Y=2184000
X5341 24 5178 ICV_13 $T=9720000 3344000 0 0 $X=9720000 $Y=3344000
X5342 24 5179 ICV_13 $T=9784000 1256000 0 0 $X=9784000 $Y=1256000
X5343 24 5180 ICV_13 $T=9928000 8680000 0 0 $X=9928000 $Y=8680000
X5344 24 5181 ICV_13 $T=10184000 2880000 0 0 $X=10184000 $Y=2880000
X5345 24 5182 ICV_13 $T=10208000 8680000 0 0 $X=10208000 $Y=8680000
X5346 24 5183 ICV_13 $T=10488000 5896000 0 0 $X=10488000 $Y=5896000
X5347 24 2353 ICV_13 $T=10808000 3808000 0 0 $X=10808000 $Y=3808000
X5348 24 5184 ICV_13 $T=10808000 4736000 0 0 $X=10808000 $Y=4736000
X5349 24 5185 ICV_13 $T=10832000 11232000 0 0 $X=10832000 $Y=11232000
X5350 24 5186 ICV_13 $T=10896000 3112000 0 0 $X=10896000 $Y=3112000
X5351 24 5187 ICV_13 $T=10912000 7984000 0 0 $X=10912000 $Y=7984000
X5352 24 5188 ICV_13 $T=11048000 6592000 0 0 $X=11048000 $Y=6592000
X5353 24 5189 ICV_13 $T=11808000 5896000 0 0 $X=11808000 $Y=5896000
X5354 24 5190 ICV_13 $T=11816000 6128000 0 0 $X=11816000 $Y=6128000
X5355 24 ICV_14 $T=1352000 5664000 1 180 $X=1168000 $Y=5664000
X5356 24 ICV_14 $T=3448000 13320000 1 180 $X=3264000 $Y=13320000
X5357 24 ICV_14 $T=5136000 8448000 1 180 $X=4952000 $Y=8448000
X5358 24 ICV_14 $T=5832000 6592000 1 180 $X=5648000 $Y=6592000
X5359 24 ICV_14 $T=10264000 7984000 1 180 $X=10080000 $Y=7984000
X5360 24 ICV_14 $T=11072000 6824000 1 180 $X=10888000 $Y=6824000
X5361 24 ICV_14 $T=11672000 2184000 1 180 $X=11488000 $Y=2184000
X5362 24 ICV_14 $T=11680000 4736000 1 180 $X=11496000 $Y=4736000
X5363 24 ICV_14 $T=11976000 2416000 1 180 $X=11792000 $Y=2416000
X5364 24 ICV_15 $T=1344000 6592000 1 180 $X=1160000 $Y=6592000
X5365 24 ICV_15 $T=2360000 7984000 1 180 $X=2176000 $Y=7984000
X5366 24 ICV_15 $T=3864000 8216000 1 180 $X=3680000 $Y=8216000
X5367 24 ICV_15 $T=5752000 5200000 1 180 $X=5568000 $Y=5200000
X5368 24 ICV_15 $T=8336000 1720000 1 180 $X=8152000 $Y=1720000
X5369 24 ICV_15 $T=8760000 6824000 1 180 $X=8576000 $Y=6824000
X5370 24 ICV_15 $T=9152000 12856000 1 180 $X=8968000 $Y=12856000
X5371 24 ICV_15 $T=10496000 6128000 1 180 $X=10312000 $Y=6128000
X5372 24 ICV_15 $T=11104000 9376000 1 180 $X=10920000 $Y=9376000
X5373 24 ICV_15 $T=11112000 7752000 1 180 $X=10928000 $Y=7752000
X5374 24 ICV_15 $T=11176000 2184000 1 180 $X=10992000 $Y=2184000
X5375 24 ICV_15 $T=11784000 9376000 1 180 $X=11600000 $Y=9376000
X5376 24 ICV_15 $T=11912000 11000000 1 180 $X=11728000 $Y=11000000
X5377 24 ICV_15 $T=11968000 8448000 1 180 $X=11784000 $Y=8448000
X5378 24 5191 ICV_16 $T=400000 5896000 0 0 $X=400000 $Y=5896000
X5379 24 5192 ICV_16 $T=464000 8216000 0 0 $X=464000 $Y=8216000
X5380 24 5193 ICV_16 $T=576000 10304000 0 0 $X=576000 $Y=10304000
X5381 24 5194 ICV_16 $T=648000 4968000 0 0 $X=648000 $Y=4968000
X5382 24 5195 ICV_16 $T=880000 4736000 0 0 $X=880000 $Y=4736000
X5383 24 5196 ICV_16 $T=952000 6360000 0 0 $X=952000 $Y=6360000
X5384 24 5197 ICV_16 $T=984000 13320000 0 0 $X=984000 $Y=13320000
X5385 24 5198 ICV_16 $T=1584000 12392000 0 0 $X=1584000 $Y=12392000
X5386 24 5199 ICV_16 $T=1864000 4040000 0 0 $X=1864000 $Y=4040000
X5387 24 5200 ICV_16 $T=1888000 3808000 0 0 $X=1888000 $Y=3808000
X5388 24 5201 ICV_16 $T=1920000 5896000 0 0 $X=1920000 $Y=5896000
X5389 24 5202 ICV_16 $T=1952000 8912000 0 0 $X=1952000 $Y=8912000
X5390 24 5203 ICV_16 $T=1968000 9144000 0 0 $X=1968000 $Y=9144000
X5391 24 5204 ICV_16 $T=1992000 8680000 0 0 $X=1992000 $Y=8680000
X5392 24 5205 ICV_16 $T=2232000 4504000 0 0 $X=2232000 $Y=4504000
X5393 24 5206 ICV_16 $T=2624000 4736000 0 0 $X=2624000 $Y=4736000
X5394 24 5207 ICV_16 $T=3048000 9840000 0 0 $X=3048000 $Y=9840000
X5395 24 5208 ICV_16 $T=3280000 9608000 0 0 $X=3280000 $Y=9608000
X5396 24 5209 ICV_16 $T=3344000 7056000 0 0 $X=3344000 $Y=7056000
X5397 24 5210 ICV_16 $T=3352000 7520000 0 0 $X=3352000 $Y=7520000
X5398 24 5211 ICV_16 $T=3440000 6360000 0 0 $X=3440000 $Y=6360000
X5399 24 5212 ICV_16 $T=3456000 2416000 0 0 $X=3456000 $Y=2416000
X5400 24 5213 ICV_16 $T=3480000 1952000 0 0 $X=3480000 $Y=1952000
X5401 24 5214 ICV_16 $T=3488000 4968000 0 0 $X=3488000 $Y=4968000
X5402 24 5215 ICV_16 $T=3488000 6128000 0 0 $X=3488000 $Y=6128000
X5403 24 5216 ICV_16 $T=3496000 5664000 0 0 $X=3496000 $Y=5664000
X5404 24 5217 ICV_16 $T=3528000 792000 0 0 $X=3528000 $Y=792000
X5405 24 5218 ICV_16 $T=3552000 4736000 0 0 $X=3552000 $Y=4736000
X5406 24 5219 ICV_16 $T=3704000 1024000 0 0 $X=3704000 $Y=1024000
X5407 24 5220 ICV_16 $T=3744000 10768000 0 0 $X=3744000 $Y=10768000
X5408 24 5221 ICV_16 $T=3760000 2184000 0 0 $X=3760000 $Y=2184000
X5409 24 5222 ICV_16 $T=3776000 7056000 0 0 $X=3776000 $Y=7056000
X5410 24 5223 ICV_16 $T=3792000 13320000 0 0 $X=3792000 $Y=13320000
X5411 24 5224 ICV_16 $T=3848000 7288000 0 0 $X=3848000 $Y=7288000
X5412 24 5225 ICV_16 $T=3960000 3344000 0 0 $X=3960000 $Y=3344000
X5413 24 5226 ICV_16 $T=4072000 11232000 0 0 $X=4072000 $Y=11232000
X5414 24 5227 ICV_16 $T=4096000 6592000 0 0 $X=4096000 $Y=6592000
X5415 24 5228 ICV_16 $T=4136000 3576000 0 0 $X=4136000 $Y=3576000
X5416 24 5229 ICV_16 $T=4472000 5664000 0 0 $X=4472000 $Y=5664000
X5417 24 5230 ICV_16 $T=4736000 9840000 0 0 $X=4736000 $Y=9840000
X5418 24 5231 ICV_16 $T=4800000 1024000 0 0 $X=4800000 $Y=1024000
X5419 24 5232 ICV_16 $T=4800000 3112000 0 0 $X=4800000 $Y=3112000
X5420 24 5233 ICV_16 $T=4808000 6360000 0 0 $X=4808000 $Y=6360000
X5421 24 5234 ICV_16 $T=4824000 560000 0 0 $X=4824000 $Y=560000
X5422 24 5235 ICV_16 $T=4880000 12856000 0 0 $X=4880000 $Y=12856000
X5423 24 5236 ICV_16 $T=4888000 6592000 0 0 $X=4888000 $Y=6592000
X5424 24 5237 ICV_16 $T=4952000 2880000 0 0 $X=4952000 $Y=2880000
X5425 24 5238 ICV_16 $T=5096000 4040000 0 0 $X=5096000 $Y=4040000
X5426 24 5239 ICV_16 $T=5112000 3344000 0 0 $X=5112000 $Y=3344000
X5427 24 5240 ICV_16 $T=5216000 4272000 0 0 $X=5216000 $Y=4272000
X5428 24 5241 ICV_16 $T=5264000 4968000 0 0 $X=5264000 $Y=4968000
X5429 24 5242 ICV_16 $T=5296000 7288000 0 0 $X=5296000 $Y=7288000
X5430 24 5243 ICV_16 $T=5352000 11464000 0 0 $X=5352000 $Y=11464000
X5431 24 5244 ICV_16 $T=5408000 12392000 0 0 $X=5408000 $Y=12392000
X5432 24 5245 ICV_16 $T=5480000 792000 0 0 $X=5480000 $Y=792000
X5433 24 5246 ICV_16 $T=5592000 7288000 0 0 $X=5592000 $Y=7288000
X5434 24 5247 ICV_16 $T=5792000 9376000 0 0 $X=5792000 $Y=9376000
X5435 24 5248 ICV_16 $T=6344000 3576000 0 0 $X=6344000 $Y=3576000
X5436 24 5249 ICV_16 $T=6344000 4736000 0 0 $X=6344000 $Y=4736000
X5437 24 2332 ICV_16 $T=6376000 4504000 0 0 $X=6376000 $Y=4504000
X5438 24 5250 ICV_16 $T=6440000 1024000 0 0 $X=6440000 $Y=1024000
X5439 24 5251 ICV_16 $T=6496000 1720000 0 0 $X=6496000 $Y=1720000
X5440 24 5252 ICV_16 $T=6504000 13088000 0 0 $X=6504000 $Y=13088000
X5441 24 5253 ICV_16 $T=6568000 13552000 0 0 $X=6568000 $Y=13552000
X5442 24 5254 ICV_16 $T=6592000 8912000 0 0 $X=6592000 $Y=8912000
X5443 24 5255 ICV_16 $T=6616000 328000 0 0 $X=6616000 $Y=328000
X5444 24 5256 ICV_16 $T=6656000 11000000 0 0 $X=6656000 $Y=11000000
X5445 24 5257 ICV_16 $T=6696000 9840000 0 0 $X=6696000 $Y=9840000
X5446 24 5258 ICV_16 $T=6704000 9608000 0 0 $X=6704000 $Y=9608000
X5447 24 5259 ICV_16 $T=6728000 792000 0 0 $X=6728000 $Y=792000
X5448 24 5260 ICV_16 $T=6752000 10768000 0 0 $X=6752000 $Y=10768000
X5449 24 5261 ICV_16 $T=6832000 7520000 0 0 $X=6832000 $Y=7520000
X5450 24 5262 ICV_16 $T=6872000 7288000 0 0 $X=6872000 $Y=7288000
X5451 24 5263 ICV_16 $T=6984000 4736000 0 0 $X=6984000 $Y=4736000
X5452 24 5264 ICV_16 $T=7096000 8448000 0 0 $X=7096000 $Y=8448000
X5453 24 5265 ICV_16 $T=7112000 12392000 0 0 $X=7112000 $Y=12392000
X5454 24 5266 ICV_16 $T=7216000 13088000 0 0 $X=7216000 $Y=13088000
X5455 24 5267 ICV_16 $T=7352000 7984000 0 0 $X=7352000 $Y=7984000
X5456 24 5268 ICV_16 $T=7408000 11696000 0 0 $X=7408000 $Y=11696000
X5457 24 5269 ICV_16 $T=7456000 5896000 0 0 $X=7456000 $Y=5896000
X5458 24 5270 ICV_16 $T=7536000 5432000 0 0 $X=7536000 $Y=5432000
X5459 24 5271 ICV_16 $T=7704000 2416000 0 0 $X=7704000 $Y=2416000
X5460 24 5272 ICV_16 $T=7760000 1952000 0 0 $X=7760000 $Y=1952000
X5461 24 5273 ICV_16 $T=7832000 792000 0 0 $X=7832000 $Y=792000
X5462 24 5274 ICV_16 $T=7880000 2648000 0 0 $X=7880000 $Y=2648000
X5463 24 5275 ICV_16 $T=7936000 12160000 0 0 $X=7936000 $Y=12160000
X5464 24 5276 ICV_16 $T=8056000 6592000 0 0 $X=8056000 $Y=6592000
X5465 24 5277 ICV_16 $T=8096000 4968000 0 0 $X=8096000 $Y=4968000
X5466 24 5278 ICV_16 $T=8096000 10768000 0 0 $X=8096000 $Y=10768000
X5467 24 5279 ICV_16 $T=8112000 11000000 0 0 $X=8112000 $Y=11000000
X5468 24 5280 ICV_16 $T=8160000 9376000 0 0 $X=8160000 $Y=9376000
X5469 24 5281 ICV_16 $T=8224000 4272000 0 0 $X=8224000 $Y=4272000
X5470 24 5282 ICV_16 $T=8240000 6824000 0 0 $X=8240000 $Y=6824000
X5471 24 5283 ICV_16 $T=8448000 8912000 0 0 $X=8448000 $Y=8912000
X5472 24 5284 ICV_16 $T=8496000 7520000 0 0 $X=8496000 $Y=7520000
X5473 24 5285 ICV_16 $T=8496000 10304000 0 0 $X=8496000 $Y=10304000
X5474 24 5286 ICV_16 $T=8656000 3344000 0 0 $X=8656000 $Y=3344000
X5475 24 5287 ICV_16 $T=8728000 3808000 0 0 $X=8728000 $Y=3808000
X5476 24 5288 ICV_16 $T=8744000 560000 0 0 $X=8744000 $Y=560000
X5477 24 5289 ICV_16 $T=8808000 4272000 0 0 $X=8808000 $Y=4272000
X5478 24 5290 ICV_16 $T=8824000 9840000 0 0 $X=8824000 $Y=9840000
X5479 24 5291 ICV_16 $T=8848000 328000 0 0 $X=8848000 $Y=328000
X5480 24 5292 ICV_16 $T=8856000 10536000 0 0 $X=8856000 $Y=10536000
X5481 24 5293 ICV_16 $T=8872000 5432000 0 0 $X=8872000 $Y=5432000
X5482 24 5294 ICV_16 $T=8904000 6360000 0 0 $X=8904000 $Y=6360000
X5483 24 4576 ICV_16 $T=8992000 5664000 0 0 $X=8992000 $Y=5664000
X5484 24 5295 ICV_16 $T=9024000 5896000 0 0 $X=9024000 $Y=5896000
X5485 24 5296 ICV_16 $T=9080000 1720000 0 0 $X=9080000 $Y=1720000
X5486 24 5297 ICV_16 $T=9160000 2184000 0 0 $X=9160000 $Y=2184000
X5487 24 5298 ICV_16 $T=9176000 8216000 0 0 $X=9176000 $Y=8216000
X5488 24 5299 ICV_16 $T=9424000 3112000 0 0 $X=9424000 $Y=3112000
X5489 24 5300 ICV_16 $T=9688000 3576000 0 0 $X=9688000 $Y=3576000
X5490 24 5301 ICV_16 $T=9744000 10304000 0 0 $X=9744000 $Y=10304000
X5491 24 5302 ICV_16 $T=9784000 10072000 0 0 $X=9784000 $Y=10072000
X5492 24 5303 ICV_16 $T=9792000 11232000 0 0 $X=9792000 $Y=11232000
X5493 24 5304 ICV_16 $T=9816000 6360000 0 0 $X=9816000 $Y=6360000
X5494 24 5305 ICV_16 $T=9896000 7520000 0 0 $X=9896000 $Y=7520000
X5495 24 5306 ICV_16 $T=9952000 11928000 0 0 $X=9952000 $Y=11928000
X5496 24 5307 ICV_16 $T=10000000 3344000 0 0 $X=10000000 $Y=3344000
X5497 24 5308 ICV_16 $T=10016000 4504000 0 0 $X=10016000 $Y=4504000
X5498 24 5309 ICV_16 $T=10088000 10072000 0 0 $X=10088000 $Y=10072000
X5499 24 5310 ICV_16 $T=10176000 3808000 0 0 $X=10176000 $Y=3808000
X5500 24 5311 ICV_16 $T=10200000 6824000 0 0 $X=10200000 $Y=6824000
X5501 24 5312 ICV_16 $T=10240000 3576000 0 0 $X=10240000 $Y=3576000
X5502 24 5313 ICV_16 $T=10448000 8216000 0 0 $X=10448000 $Y=8216000
X5503 24 5314 ICV_16 $T=10480000 13320000 0 0 $X=10480000 $Y=13320000
X5504 24 5315 ICV_16 $T=10520000 5200000 0 0 $X=10520000 $Y=5200000
X5505 24 5316 ICV_16 $T=10576000 5432000 0 0 $X=10576000 $Y=5432000
X5506 24 5317 ICV_16 $T=10584000 2184000 0 0 $X=10584000 $Y=2184000
X5507 24 5318 ICV_16 $T=10696000 7520000 0 0 $X=10696000 $Y=7520000
X5508 24 5319 ICV_16 $T=11216000 12392000 0 0 $X=11216000 $Y=12392000
X5509 24 5320 ICV_16 $T=11288000 2648000 0 0 $X=11288000 $Y=2648000
X5510 24 5321 ICV_16 $T=11288000 11696000 0 0 $X=11288000 $Y=11696000
X5511 24 5322 ICV_16 $T=11616000 4272000 0 0 $X=11616000 $Y=4272000
X5512 24 5323 ICV_16 $T=11744000 3808000 0 0 $X=11744000 $Y=3808000
X5513 24 2588 ICV_17 $T=1944000 13320000 0 0 $X=1944000 $Y=13320000
X5514 24 3067 ICV_17 $T=2416000 9144000 0 0 $X=2416000 $Y=9144000
X5515 24 5324 ICV_17 $T=2592000 7056000 0 0 $X=2592000 $Y=7056000
X5516 24 5325 ICV_17 $T=4296000 1256000 0 0 $X=4296000 $Y=1256000
X5517 24 464 ICV_17 $T=4368000 8680000 0 0 $X=4368000 $Y=8680000
X5518 24 5051 ICV_17 $T=4520000 5200000 0 0 $X=4520000 $Y=5200000
X5519 24 3201 ICV_17 $T=4592000 12624000 0 0 $X=4592000 $Y=12624000
X5520 24 510 ICV_17 $T=5048000 96000 0 0 $X=5048000 $Y=96000
X5521 24 3846 ICV_17 $T=5256000 5896000 0 0 $X=5256000 $Y=5896000
X5522 24 2332 ICV_17 $T=5824000 4504000 0 0 $X=5824000 $Y=4504000
X5523 24 2333 ICV_17 $T=6032000 7056000 0 0 $X=6032000 $Y=7056000
X5524 24 5326 ICV_17 $T=6040000 1952000 0 0 $X=6040000 $Y=1952000
X5525 24 5327 ICV_17 $T=6912000 7056000 0 0 $X=6912000 $Y=7056000
X5526 24 744 ICV_17 $T=7664000 8216000 0 0 $X=7664000 $Y=8216000
X5527 24 4013 ICV_17 $T=9224000 4272000 0 0 $X=9224000 $Y=4272000
X5528 24 1907 ICV_17 $T=9328000 4736000 0 0 $X=9328000 $Y=4736000
X5529 24 3542 ICV_17 $T=9936000 1952000 0 0 $X=9936000 $Y=1952000
X5530 24 27 ICV_17 $T=10120000 328000 0 0 $X=10120000 $Y=328000
X5531 24 5328 ICV_17 $T=10344000 3112000 0 0 $X=10344000 $Y=3112000
X5532 24 5329 ICV_17 $T=10592000 13552000 0 0 $X=10592000 $Y=13552000
X5533 24 2883 ICV_17 $T=10744000 12392000 0 0 $X=10744000 $Y=12392000
X5534 24 2062 ICV_17 $T=10856000 8448000 0 0 $X=10856000 $Y=8448000
X5535 24 3658 ICV_17 $T=11616000 3112000 0 0 $X=11616000 $Y=3112000
X5536 24 4094 ICV_17 $T=11728000 6360000 0 0 $X=11728000 $Y=6360000
X5537 24 5330 xnor2 $T=279000 3576000 1 180 $X=216000 $Y=3576000
X5538 24 5331 xnor2 $T=279000 4040000 1 180 $X=216000 $Y=4040000
X5539 24 5332 xnor2 $T=375000 2184000 1 180 $X=312000 $Y=2184000
X5540 24 5333 xnor2 $T=384000 3808000 0 0 $X=384000 $Y=3808000
X5541 24 5334 xnor2 $T=503000 3576000 1 180 $X=440000 $Y=3576000
X5542 24 5335 xnor2 $T=568000 96000 0 0 $X=568000 $Y=96000
X5543 24 5336 xnor2 $T=631000 3808000 1 180 $X=568000 $Y=3808000
X5544 24 5337 xnor2 $T=679000 2184000 1 180 $X=616000 $Y=2184000
X5545 24 5338 xnor2 $T=695000 1024000 1 180 $X=632000 $Y=1024000
X5546 24 5339 xnor2 $T=704000 2416000 0 0 $X=704000 $Y=2416000
X5547 24 5340 xnor2 $T=823000 328000 1 180 $X=760000 $Y=328000
X5548 24 5341 xnor2 $T=776000 3112000 0 0 $X=776000 $Y=3112000
X5549 24 5342 xnor2 $T=776000 4272000 0 0 $X=776000 $Y=4272000
X5550 24 5343 xnor2 $T=792000 2880000 0 0 $X=792000 $Y=2880000
X5551 24 5344 xnor2 $T=1103000 2648000 1 180 $X=1040000 $Y=2648000
X5552 24 5345 xnor2 $T=1184000 2184000 0 0 $X=1184000 $Y=2184000
X5553 24 5346 xnor2 $T=1192000 2880000 0 0 $X=1192000 $Y=2880000
X5554 24 5347 xnor2 $T=1240000 2648000 0 0 $X=1240000 $Y=2648000
X5555 24 5348 xnor2 $T=1367000 2648000 1 180 $X=1304000 $Y=2648000
X5556 24 5349 xnor2 $T=1320000 3808000 0 0 $X=1320000 $Y=3808000
X5557 24 5350 xnor2 $T=1431000 2184000 1 180 $X=1368000 $Y=2184000
X5558 24 5351 xnor2 $T=1447000 3808000 1 180 $X=1384000 $Y=3808000
X5559 24 5352 xnor2 $T=1400000 1256000 0 0 $X=1400000 $Y=1256000
X5560 24 5353 xnor2 $T=1472000 792000 0 0 $X=1472000 $Y=792000
X5561 24 5354 xnor2 $T=1512000 2880000 0 0 $X=1512000 $Y=2880000
X5562 24 5355 xnor2 $T=1895000 1256000 1 180 $X=1832000 $Y=1256000
X5563 24 5356 xnor2 $T=1936000 328000 0 0 $X=1936000 $Y=328000
X5564 24 5357 xnor2 $T=2143000 1256000 1 180 $X=2080000 $Y=1256000
X5565 24 5358 xnor2 $T=2216000 1488000 0 0 $X=2216000 $Y=1488000
X5566 24 5359 xnor2 $T=2344000 328000 0 0 $X=2344000 $Y=328000
X5567 24 5360 xnor2 $T=2623000 2184000 1 180 $X=2560000 $Y=2184000
X5568 24 5361 xnor2 $T=2631000 1488000 1 180 $X=2568000 $Y=1488000
X5569 24 5362 xnor2 $T=2703000 96000 1 180 $X=2640000 $Y=96000
X5570 24 5363 xnor2 $T=2831000 1720000 1 180 $X=2768000 $Y=1720000
X5571 24 5364 xnor2 $T=2816000 2416000 0 0 $X=2816000 $Y=2416000
X5572 24 5365 xnor2 $T=2911000 1256000 1 180 $X=2848000 $Y=1256000
X5573 24 5366 xnor2 $T=2960000 792000 0 0 $X=2960000 $Y=792000
X5574 24 5367 xnor2 $T=3056000 792000 0 0 $X=3056000 $Y=792000
X5575 24 5368 xnor2 $T=3056000 1720000 0 0 $X=3056000 $Y=1720000
X5576 24 5369 xnor2 $T=3072000 1256000 0 0 $X=3072000 $Y=1256000
X5577 24 5370 xnor2 $T=3552000 328000 0 0 $X=3552000 $Y=328000
X5578 24 5371 xnor2 $T=3640000 96000 0 0 $X=3640000 $Y=96000
X5579 24 5372 xnor2 $T=3704000 328000 0 0 $X=3704000 $Y=328000
X5580 24 5373 xnor2 $T=4080000 96000 0 0 $X=4080000 $Y=96000
X5581 24 5374 xnor2 $T=10711000 1024000 1 180 $X=10648000 $Y=1024000
X5582 24 5375 xnor2 $T=10839000 792000 1 180 $X=10776000 $Y=792000
X5583 24 5376 xnor2 $T=10936000 560000 0 0 $X=10936000 $Y=560000
X5584 24 5377 xnor2 $T=11720000 7056000 0 0 $X=11720000 $Y=7056000
X5585 24 5378 ICV_18 $T=376000 792000 0 0 $X=376000 $Y=792000
X5586 24 5379 ICV_18 $T=784000 2416000 0 0 $X=784000 $Y=2416000
X5587 24 5380 ICV_18 $T=800000 3576000 0 0 $X=800000 $Y=3576000
X5588 24 5381 ICV_18 $T=816000 4040000 0 0 $X=816000 $Y=4040000
X5589 24 5382 ICV_18 $T=1072000 560000 0 0 $X=1072000 $Y=560000
X5590 24 5383 ICV_18 $T=2160000 792000 0 0 $X=2160000 $Y=792000
X5591 24 5384 ICV_18 $T=2208000 560000 0 0 $X=2208000 $Y=560000
X5592 24 5385 ICV_18 $T=2384000 1024000 0 0 $X=2384000 $Y=1024000
X5593 24 5386 ICV_18 $T=3128000 96000 0 0 $X=3128000 $Y=96000
X5594 24 5387 ICV_18 $T=3792000 96000 0 0 $X=3792000 $Y=96000
X5595 24 5388 ICV_18 $T=4232000 96000 0 0 $X=4232000 $Y=96000
X5596 24 2356 ICV_18 $T=11488000 3112000 0 0 $X=11488000 $Y=3112000
X5597 24 5389 ICV_18 $T=11704000 6824000 0 0 $X=11704000 $Y=6824000
X5598 24 xor2 $T=152000 3808000 0 0 $X=152000 $Y=3808000
X5599 24 xor2 $T=256000 3808000 0 0 $X=256000 $Y=3808000
X5600 24 xor2 $T=440000 3344000 0 0 $X=440000 $Y=3344000
X5601 24 xor2 $T=632000 96000 0 0 $X=632000 $Y=96000
X5602 24 xor2 $T=910000 3112000 1 180 $X=840000 $Y=3112000
X5603 24 xor2 $T=912000 560000 0 0 $X=912000 $Y=560000
X5604 24 xor2 $T=982000 3112000 1 180 $X=912000 $Y=3112000
X5605 24 xor2 $T=1054000 3112000 1 180 $X=984000 $Y=3112000
X5606 24 xor2 $T=1142000 2880000 1 180 $X=1072000 $Y=2880000
X5607 24 xor2 $T=1240000 1256000 0 0 $X=1240000 $Y=1256000
X5608 24 xor2 $T=1326000 2880000 1 180 $X=1256000 $Y=2880000
X5609 24 xor2 $T=1334000 5200000 1 180 $X=1264000 $Y=5200000
X5610 24 xor2 $T=1376000 3112000 0 0 $X=1376000 $Y=3112000
X5611 24 xor2 $T=1454000 4040000 1 180 $X=1384000 $Y=4040000
X5612 24 xor2 $T=1614000 1720000 1 180 $X=1544000 $Y=1720000
X5613 24 xor2 $T=2280000 96000 0 0 $X=2280000 $Y=96000
X5614 24 xor2 $T=2694000 560000 1 180 $X=2624000 $Y=560000
X5615 24 xor2 $T=2774000 96000 1 180 $X=2704000 $Y=96000
X5616 24 xor2 $T=2712000 2416000 0 0 $X=2712000 $Y=2416000
X5617 24 xor2 $T=2846000 2184000 1 180 $X=2776000 $Y=2184000
X5618 24 xor2 $T=2776000 2648000 0 0 $X=2776000 $Y=2648000
X5619 24 xor2 $T=2982000 1256000 1 180 $X=2912000 $Y=1256000
X5620 24 xor2 $T=2952000 1720000 0 0 $X=2952000 $Y=1720000
X5621 24 xor2 $T=3038000 96000 1 180 $X=2968000 $Y=96000
X5622 24 xor2 $T=3070000 1488000 1 180 $X=3000000 $Y=1488000
X5623 24 xor2 $T=3416000 96000 0 0 $X=3416000 $Y=96000
X5624 24 xor2 $T=4206000 328000 1 180 $X=4136000 $Y=328000
X5625 24 xor2 $T=10632000 792000 0 0 $X=10632000 $Y=792000
X5626 24 xor2 $T=10704000 792000 0 0 $X=10704000 $Y=792000
X5627 24 xor2 $T=11014000 328000 1 180 $X=10944000 $Y=328000
X5628 24 xor2 $T=11488000 6592000 0 0 $X=11488000 $Y=6592000
X5629 24 xor2 $T=11646000 1720000 1 180 $X=11576000 $Y=1720000
X5630 24 xor2 $T=11616000 6592000 0 0 $X=11616000 $Y=6592000
X5631 24 5390 ICV_19 $T=152000 4736000 0 0 $X=152000 $Y=4736000
X5632 24 5391 ICV_19 $T=152000 4968000 0 0 $X=152000 $Y=4968000
X5633 24 5392 ICV_19 $T=152000 5896000 0 0 $X=152000 $Y=5896000
X5634 24 5393 ICV_19 $T=152000 6128000 0 0 $X=152000 $Y=6128000
X5635 24 5394 ICV_19 $T=152000 6592000 0 0 $X=152000 $Y=6592000
X5636 24 5395 ICV_19 $T=152000 6824000 0 0 $X=152000 $Y=6824000
X5637 24 5396 ICV_19 $T=152000 7056000 0 0 $X=152000 $Y=7056000
X5638 24 5397 ICV_19 $T=152000 7520000 0 0 $X=152000 $Y=7520000
X5639 24 5398 ICV_19 $T=152000 7984000 0 0 $X=152000 $Y=7984000
X5640 24 5399 ICV_19 $T=152000 8216000 0 0 $X=152000 $Y=8216000
X5641 24 5400 ICV_19 $T=152000 8448000 0 0 $X=152000 $Y=8448000
X5642 24 5401 ICV_19 $T=152000 11464000 0 0 $X=152000 $Y=11464000
X5643 24 5402 ICV_19 $T=152000 12392000 0 0 $X=152000 $Y=12392000
X5644 24 5403 ICV_19 $T=152000 12856000 0 0 $X=152000 $Y=12856000
X5645 24 5404 ICV_19 $T=152000 13320000 0 0 $X=152000 $Y=13320000
X5646 24 5405 ICV_19 $T=192000 8912000 0 0 $X=192000 $Y=8912000
X5647 24 5406 ICV_19 $T=216000 4504000 0 0 $X=216000 $Y=4504000
X5648 24 5407 ICV_19 $T=216000 10304000 0 0 $X=216000 $Y=10304000
X5649 24 5408 ICV_19 $T=216000 13088000 0 0 $X=216000 $Y=13088000
X5650 24 5409 ICV_19 $T=232000 12160000 0 0 $X=232000 $Y=12160000
X5651 24 5410 ICV_19 $T=400000 6592000 0 0 $X=400000 $Y=6592000
X5652 24 5411 ICV_19 $T=400000 7984000 0 0 $X=400000 $Y=7984000
X5653 24 5412 ICV_19 $T=400000 11000000 0 0 $X=400000 $Y=11000000
X5654 24 5413 ICV_19 $T=400000 12856000 0 0 $X=400000 $Y=12856000
X5655 24 5414 ICV_19 $T=424000 11928000 0 0 $X=424000 $Y=11928000
X5656 24 5415 ICV_19 $T=432000 6360000 0 0 $X=432000 $Y=6360000
X5657 24 5416 ICV_19 $T=440000 8912000 0 0 $X=440000 $Y=8912000
X5658 24 5417 ICV_19 $T=464000 7056000 0 0 $X=464000 $Y=7056000
X5659 24 5418 ICV_19 $T=512000 13088000 0 0 $X=512000 $Y=13088000
X5660 24 5419 ICV_19 $T=616000 5200000 0 0 $X=616000 $Y=5200000
X5661 24 5420 ICV_19 $T=624000 10536000 0 0 $X=624000 $Y=10536000
X5662 24 5421 ICV_19 $T=744000 5664000 0 0 $X=744000 $Y=5664000
X5663 24 5422 ICV_19 $T=808000 4504000 0 0 $X=808000 $Y=4504000
X5664 24 5423 ICV_19 $T=832000 7520000 0 0 $X=832000 $Y=7520000
X5665 24 5424 ICV_19 $T=840000 7056000 0 0 $X=840000 $Y=7056000
X5666 24 5425 ICV_19 $T=856000 6592000 0 0 $X=856000 $Y=6592000
X5667 24 5426 ICV_19 $T=856000 7984000 0 0 $X=856000 $Y=7984000
X5668 24 5427 ICV_19 $T=872000 10536000 0 0 $X=872000 $Y=10536000
X5669 24 5428 ICV_19 $T=888000 8448000 0 0 $X=888000 $Y=8448000
X5670 24 5429 ICV_19 $T=904000 11000000 0 0 $X=904000 $Y=11000000
X5671 24 5430 ICV_19 $T=928000 9608000 0 0 $X=928000 $Y=9608000
X5672 24 5431 ICV_19 $T=928000 11464000 0 0 $X=928000 $Y=11464000
X5673 24 5432 ICV_19 $T=936000 8912000 0 0 $X=936000 $Y=8912000
X5674 24 5433 ICV_19 $T=968000 7752000 0 0 $X=968000 $Y=7752000
X5675 24 5434 ICV_19 $T=1088000 8680000 0 0 $X=1088000 $Y=8680000
X5676 24 5435 ICV_19 $T=1152000 9840000 0 0 $X=1152000 $Y=9840000
X5677 24 5436 ICV_19 $T=1216000 12392000 0 0 $X=1216000 $Y=12392000
X5678 24 5437 ICV_19 $T=1384000 12624000 0 0 $X=1384000 $Y=12624000
X5679 24 5438 ICV_19 $T=1528000 4968000 0 0 $X=1528000 $Y=4968000
X5680 24 5439 ICV_19 $T=1536000 9376000 0 0 $X=1536000 $Y=9376000
X5681 24 5440 ICV_19 $T=1584000 12160000 0 0 $X=1584000 $Y=12160000
X5682 24 5441 ICV_19 $T=1616000 10768000 0 0 $X=1616000 $Y=10768000
X5683 24 5442 ICV_19 $T=1640000 8912000 0 0 $X=1640000 $Y=8912000
X5684 24 5443 ICV_19 $T=1648000 8680000 0 0 $X=1648000 $Y=8680000
X5685 24 5444 ICV_19 $T=1656000 9144000 0 0 $X=1656000 $Y=9144000
X5686 24 5445 ICV_19 $T=1960000 4272000 0 0 $X=1960000 $Y=4272000
X5687 24 5446 ICV_19 $T=2032000 10536000 0 0 $X=2032000 $Y=10536000
X5688 24 5447 ICV_19 $T=2048000 11928000 0 0 $X=2048000 $Y=11928000
X5689 24 5448 ICV_19 $T=2088000 5200000 0 0 $X=2088000 $Y=5200000
X5690 24 5449 ICV_19 $T=2120000 9376000 0 0 $X=2120000 $Y=9376000
X5691 24 5450 ICV_19 $T=2144000 13552000 0 0 $X=2144000 $Y=13552000
X5692 24 5451 ICV_19 $T=2152000 4736000 0 0 $X=2152000 $Y=4736000
X5693 24 5452 ICV_19 $T=2192000 12856000 0 0 $X=2192000 $Y=12856000
X5694 24 5453 ICV_19 $T=2248000 9608000 0 0 $X=2248000 $Y=9608000
X5695 24 5454 ICV_19 $T=2264000 11696000 0 0 $X=2264000 $Y=11696000
X5696 24 5455 ICV_19 $T=2280000 7056000 0 0 $X=2280000 $Y=7056000
X5697 24 5456 ICV_19 $T=2296000 7520000 0 0 $X=2296000 $Y=7520000
X5698 24 5457 ICV_19 $T=2336000 5200000 0 0 $X=2336000 $Y=5200000
X5699 24 5458 ICV_19 $T=2448000 3344000 0 0 $X=2448000 $Y=3344000
X5700 24 5459 ICV_19 $T=2448000 6360000 0 0 $X=2448000 $Y=6360000
X5701 24 5460 ICV_19 $T=2448000 12392000 0 0 $X=2448000 $Y=12392000
X5702 24 5461 ICV_19 $T=2464000 6824000 0 0 $X=2464000 $Y=6824000
X5703 24 5462 ICV_19 $T=2488000 8680000 0 0 $X=2488000 $Y=8680000
X5704 24 5463 ICV_19 $T=2560000 8912000 0 0 $X=2560000 $Y=8912000
X5705 24 5464 ICV_19 $T=2576000 7520000 0 0 $X=2576000 $Y=7520000
X5706 24 5465 ICV_19 $T=2576000 8448000 0 0 $X=2576000 $Y=8448000
X5707 24 5466 ICV_19 $T=2736000 12392000 0 0 $X=2736000 $Y=12392000
X5708 24 5467 ICV_19 $T=2792000 10072000 0 0 $X=2792000 $Y=10072000
X5709 24 5468 ICV_19 $T=2864000 4968000 0 0 $X=2864000 $Y=4968000
X5710 24 5469 ICV_19 $T=2864000 5200000 0 0 $X=2864000 $Y=5200000
X5711 24 5470 ICV_19 $T=2896000 6592000 0 0 $X=2896000 $Y=6592000
X5712 24 5324 ICV_19 $T=2960000 7056000 0 0 $X=2960000 $Y=7056000
X5713 24 5471 ICV_19 $T=3008000 6824000 0 0 $X=3008000 $Y=6824000
X5714 24 5472 ICV_19 $T=3104000 7520000 0 0 $X=3104000 $Y=7520000
X5715 24 5473 ICV_19 $T=3120000 1720000 0 0 $X=3120000 $Y=1720000
X5716 24 5474 ICV_19 $T=3136000 1256000 0 0 $X=3136000 $Y=1256000
X5717 24 5475 ICV_19 $T=3144000 2416000 0 0 $X=3144000 $Y=2416000
X5718 24 5476 ICV_19 $T=3144000 6592000 0 0 $X=3144000 $Y=6592000
X5719 24 5477 ICV_19 $T=3152000 7752000 0 0 $X=3152000 $Y=7752000
X5720 24 5478 ICV_19 $T=3168000 1952000 0 0 $X=3168000 $Y=1952000
X5721 24 5479 ICV_19 $T=3176000 11232000 0 0 $X=3176000 $Y=11232000
X5722 24 5480 ICV_19 $T=3184000 8216000 0 0 $X=3184000 $Y=8216000
X5723 24 5481 ICV_19 $T=3192000 1488000 0 0 $X=3192000 $Y=1488000
X5724 24 5482 ICV_19 $T=3200000 2184000 0 0 $X=3200000 $Y=2184000
X5725 24 5483 ICV_19 $T=3216000 8448000 0 0 $X=3216000 $Y=8448000
X5726 24 5484 ICV_19 $T=3304000 4736000 0 0 $X=3304000 $Y=4736000
X5727 24 5485 ICV_19 $T=3320000 9840000 0 0 $X=3320000 $Y=9840000
X5728 24 5486 ICV_19 $T=3400000 7752000 0 0 $X=3400000 $Y=7752000
X5729 24 5487 ICV_19 $T=3424000 5200000 0 0 $X=3424000 $Y=5200000
X5730 24 5488 ICV_19 $T=3440000 1488000 0 0 $X=3440000 $Y=1488000
X5731 24 5489 ICV_19 $T=3440000 11928000 0 0 $X=3440000 $Y=11928000
X5732 24 5490 ICV_19 $T=3464000 11696000 0 0 $X=3464000 $Y=11696000
X5733 24 5491 ICV_19 $T=3480000 7288000 0 0 $X=3480000 $Y=7288000
X5734 24 5492 ICV_19 $T=3624000 8680000 0 0 $X=3624000 $Y=8680000
X5735 24 5493 ICV_19 $T=3648000 3344000 0 0 $X=3648000 $Y=3344000
X5736 24 5494 ICV_19 $T=3696000 560000 0 0 $X=3696000 $Y=560000
X5737 24 5495 ICV_19 $T=3760000 13552000 0 0 $X=3760000 $Y=13552000
X5738 24 5496 ICV_19 $T=3776000 12160000 0 0 $X=3776000 $Y=12160000
X5739 24 5497 ICV_19 $T=3800000 12624000 0 0 $X=3800000 $Y=12624000
X5740 24 5498 ICV_19 $T=4000000 9840000 0 0 $X=4000000 $Y=9840000
X5741 24 5499 ICV_19 $T=4016000 9376000 0 0 $X=4016000 $Y=9376000
X5742 24 5500 ICV_19 $T=4040000 5664000 0 0 $X=4040000 $Y=5664000
X5743 24 5501 ICV_19 $T=4072000 9144000 0 0 $X=4072000 $Y=9144000
X5744 24 5502 ICV_19 $T=4088000 2416000 0 0 $X=4088000 $Y=2416000
X5745 24 5503 ICV_19 $T=4096000 4968000 0 0 $X=4096000 $Y=4968000
X5746 24 5504 ICV_19 $T=4136000 6128000 0 0 $X=4136000 $Y=6128000
X5747 24 5505 ICV_19 $T=4152000 5432000 0 0 $X=4152000 $Y=5432000
X5748 24 5506 ICV_19 $T=4176000 2648000 0 0 $X=4176000 $Y=2648000
X5749 24 5507 ICV_19 $T=4216000 4504000 0 0 $X=4216000 $Y=4504000
X5750 24 5508 ICV_19 $T=4416000 7520000 0 0 $X=4416000 $Y=7520000
X5751 24 5509 ICV_19 $T=4504000 5896000 0 0 $X=4504000 $Y=5896000
X5752 24 5510 ICV_19 $T=4504000 12392000 0 0 $X=4504000 $Y=12392000
X5753 24 5511 ICV_19 $T=4728000 9376000 0 0 $X=4728000 $Y=9376000
X5754 24 5512 ICV_19 $T=4760000 10304000 0 0 $X=4760000 $Y=10304000
X5755 24 5513 ICV_19 $T=4776000 10768000 0 0 $X=4776000 $Y=10768000
X5756 24 5514 ICV_19 $T=4800000 792000 0 0 $X=4800000 $Y=792000
X5757 24 5515 ICV_19 $T=4816000 1720000 0 0 $X=4816000 $Y=1720000
X5758 24 5516 ICV_19 $T=4832000 10536000 0 0 $X=4832000 $Y=10536000
X5759 24 5517 ICV_19 $T=4856000 11696000 0 0 $X=4856000 $Y=11696000
X5760 24 5518 ICV_19 $T=4872000 7984000 0 0 $X=4872000 $Y=7984000
X5761 24 5519 ICV_19 $T=4936000 11928000 0 0 $X=4936000 $Y=11928000
X5762 24 5520 ICV_19 $T=5040000 3112000 0 0 $X=5040000 $Y=3112000
X5763 24 5521 ICV_19 $T=5064000 9376000 0 0 $X=5064000 $Y=9376000
X5764 24 5522 ICV_19 $T=5120000 7984000 0 0 $X=5120000 $Y=7984000
X5765 24 5523 ICV_19 $T=5184000 7752000 0 0 $X=5184000 $Y=7752000
X5766 24 5524 ICV_19 $T=5240000 3576000 0 0 $X=5240000 $Y=3576000
X5767 24 5525 ICV_19 $T=5352000 10768000 0 0 $X=5352000 $Y=10768000
X5768 24 5526 ICV_19 $T=5360000 11232000 0 0 $X=5360000 $Y=11232000
X5769 24 5527 ICV_19 $T=5504000 328000 0 0 $X=5504000 $Y=328000
X5770 24 5528 ICV_19 $T=5592000 11464000 0 0 $X=5592000 $Y=11464000
X5771 24 5529 ICV_19 $T=5624000 11696000 0 0 $X=5624000 $Y=11696000
X5772 24 5530 ICV_19 $T=5632000 2416000 0 0 $X=5632000 $Y=2416000
X5773 24 5531 ICV_19 $T=5640000 2880000 0 0 $X=5640000 $Y=2880000
X5774 24 5532 ICV_19 $T=5840000 10536000 0 0 $X=5840000 $Y=10536000
X5775 24 5533 ICV_19 $T=5936000 1720000 0 0 $X=5936000 $Y=1720000
X5776 24 5534 ICV_19 $T=6184000 1720000 0 0 $X=6184000 $Y=1720000
X5777 24 5535 ICV_19 $T=6248000 328000 0 0 $X=6248000 $Y=328000
X5778 24 5536 ICV_19 $T=6344000 2880000 0 0 $X=6344000 $Y=2880000
X5779 24 5537 ICV_19 $T=6344000 11232000 0 0 $X=6344000 $Y=11232000
X5780 24 5538 ICV_19 $T=6384000 6592000 0 0 $X=6384000 $Y=6592000
X5781 24 5539 ICV_19 $T=6384000 9840000 0 0 $X=6384000 $Y=9840000
X5782 24 5540 ICV_19 $T=6416000 560000 0 0 $X=6416000 $Y=560000
X5783 24 5541 ICV_19 $T=6416000 10768000 0 0 $X=6416000 $Y=10768000
X5784 24 5542 ICV_19 $T=6440000 9144000 0 0 $X=6440000 $Y=9144000
X5785 24 5543 ICV_19 $T=6448000 10072000 0 0 $X=6448000 $Y=10072000
X5786 24 5544 ICV_19 $T=6464000 3112000 0 0 $X=6464000 $Y=3112000
X5787 24 5545 ICV_19 $T=6504000 9376000 0 0 $X=6504000 $Y=9376000
X5788 24 5546 ICV_19 $T=6528000 12160000 0 0 $X=6528000 $Y=12160000
X5789 24 5547 ICV_19 $T=6536000 12392000 0 0 $X=6536000 $Y=12392000
X5790 24 5548 ICV_19 $T=6632000 12856000 0 0 $X=6632000 $Y=12856000
X5791 24 5549 ICV_19 $T=6632000 13320000 0 0 $X=6632000 $Y=13320000
X5792 24 5550 ICV_19 $T=6672000 1488000 0 0 $X=6672000 $Y=1488000
X5793 24 5551 ICV_19 $T=6688000 9144000 0 0 $X=6688000 $Y=9144000
X5794 24 5552 ICV_19 $T=6832000 10536000 0 0 $X=6832000 $Y=10536000
X5795 24 5553 ICV_19 $T=6952000 10304000 0 0 $X=6952000 $Y=10304000
X5796 24 5554 ICV_19 $T=7144000 5664000 0 0 $X=7144000 $Y=5664000
X5797 24 5555 ICV_19 $T=7176000 6824000 0 0 $X=7176000 $Y=6824000
X5798 24 5556 ICV_19 $T=7392000 2416000 0 0 $X=7392000 $Y=2416000
X5799 24 5557 ICV_19 $T=7680000 6824000 0 0 $X=7680000 $Y=6824000
X5800 24 5558 ICV_19 $T=7720000 7056000 0 0 $X=7720000 $Y=7056000
X5801 24 5559 ICV_19 $T=7728000 2184000 0 0 $X=7728000 $Y=2184000
X5802 24 5560 ICV_19 $T=7784000 4968000 0 0 $X=7784000 $Y=4968000
X5803 24 5561 ICV_19 $T=7840000 13552000 0 0 $X=7840000 $Y=13552000
X5804 24 5562 ICV_19 $T=7848000 5664000 0 0 $X=7848000 $Y=5664000
X5805 24 5563 ICV_19 $T=7872000 10536000 0 0 $X=7872000 $Y=10536000
X5806 24 5564 ICV_19 $T=7880000 10304000 0 0 $X=7880000 $Y=10304000
X5807 24 5565 ICV_19 $T=7912000 3112000 0 0 $X=7912000 $Y=3112000
X5808 24 5566 ICV_19 $T=7912000 4272000 0 0 $X=7912000 $Y=4272000
X5809 24 5567 ICV_19 $T=7912000 9840000 0 0 $X=7912000 $Y=9840000
X5810 24 5568 ICV_19 $T=7928000 6824000 0 0 $X=7928000 $Y=6824000
X5811 24 5569 ICV_19 $T=7968000 9144000 0 0 $X=7968000 $Y=9144000
X5812 24 5570 ICV_19 $T=7976000 9608000 0 0 $X=7976000 $Y=9608000
X5813 24 5571 ICV_19 $T=8008000 8448000 0 0 $X=8008000 $Y=8448000
X5814 24 5572 ICV_19 $T=8016000 13320000 0 0 $X=8016000 $Y=13320000
X5815 24 5573 ICV_19 $T=8024000 8680000 0 0 $X=8024000 $Y=8680000
X5816 24 5574 ICV_19 $T=8072000 10072000 0 0 $X=8072000 $Y=10072000
X5817 24 5575 ICV_19 $T=8080000 8912000 0 0 $X=8080000 $Y=8912000
X5818 24 5576 ICV_19 $T=8128000 13552000 0 0 $X=8128000 $Y=13552000
X5819 24 5577 ICV_19 $T=8160000 8216000 0 0 $X=8160000 $Y=8216000
X5820 24 5578 ICV_19 $T=8224000 9608000 0 0 $X=8224000 $Y=9608000
X5821 24 5579 ICV_19 $T=8232000 13088000 0 0 $X=8232000 $Y=13088000
X5822 24 5580 ICV_19 $T=8280000 9144000 0 0 $X=8280000 $Y=9144000
X5823 24 5581 ICV_19 $T=8344000 3344000 0 0 $X=8344000 $Y=3344000
X5824 24 5582 ICV_19 $T=8528000 7056000 0 0 $X=8528000 $Y=7056000
X5825 24 5583 ICV_19 $T=8528000 9144000 0 0 $X=8528000 $Y=9144000
X5826 24 5584 ICV_19 $T=8544000 11696000 0 0 $X=8544000 $Y=11696000
X5827 24 5585 ICV_19 $T=8608000 7288000 0 0 $X=8608000 $Y=7288000
X5828 24 5586 ICV_19 $T=8624000 11928000 0 0 $X=8624000 $Y=11928000
X5829 24 5587 ICV_19 $T=8688000 6128000 0 0 $X=8688000 $Y=6128000
X5830 24 5588 ICV_19 $T=8712000 5896000 0 0 $X=8712000 $Y=5896000
X5831 24 5589 ICV_19 $T=8744000 4040000 0 0 $X=8744000 $Y=4040000
X5832 24 5590 ICV_19 $T=8808000 8680000 0 0 $X=8808000 $Y=8680000
X5833 24 5591 ICV_19 $T=8816000 8912000 0 0 $X=8816000 $Y=8912000
X5834 24 5592 ICV_19 $T=8864000 7056000 0 0 $X=8864000 $Y=7056000
X5835 24 5593 ICV_19 $T=8928000 7984000 0 0 $X=8928000 $Y=7984000
X5836 24 5594 ICV_19 $T=9016000 7288000 0 0 $X=9016000 $Y=7288000
X5837 24 5595 ICV_19 $T=9368000 4504000 0 0 $X=9368000 $Y=4504000
X5838 24 5596 ICV_19 $T=9368000 9144000 0 0 $X=9368000 $Y=9144000
X5839 24 5597 ICV_19 $T=9448000 11928000 0 0 $X=9448000 $Y=11928000
X5840 24 5598 ICV_19 $T=9472000 8216000 0 0 $X=9472000 $Y=8216000
X5841 24 5599 ICV_19 $T=9472000 10072000 0 0 $X=9472000 $Y=10072000
X5842 24 5600 ICV_19 $T=9544000 11464000 0 0 $X=9544000 $Y=11464000
X5843 24 5601 ICV_19 $T=9568000 7056000 0 0 $X=9568000 $Y=7056000
X5844 24 5602 ICV_19 $T=9576000 5896000 0 0 $X=9576000 $Y=5896000
X5845 24 5603 ICV_19 $T=9616000 8448000 0 0 $X=9616000 $Y=8448000
X5846 24 5604 ICV_19 $T=9680000 11000000 0 0 $X=9680000 $Y=11000000
X5847 24 5605 ICV_19 $T=9712000 12392000 0 0 $X=9712000 $Y=12392000
X5848 24 5606 ICV_19 $T=9728000 1024000 0 0 $X=9728000 $Y=1024000
X5849 24 5607 ICV_19 $T=9760000 9144000 0 0 $X=9760000 $Y=9144000
X5850 24 5608 ICV_19 $T=9776000 7984000 0 0 $X=9776000 $Y=7984000
X5851 24 5609 ICV_19 $T=9792000 9608000 0 0 $X=9792000 $Y=9608000
X5852 24 5610 ICV_19 $T=9840000 13320000 0 0 $X=9840000 $Y=13320000
X5853 24 5611 ICV_19 $T=9848000 13552000 0 0 $X=9848000 $Y=13552000
X5854 24 5612 ICV_19 $T=10032000 11232000 0 0 $X=10032000 $Y=11232000
X5855 24 5613 ICV_19 $T=10048000 11696000 0 0 $X=10048000 $Y=11696000
X5856 24 5614 ICV_19 $T=10096000 13552000 0 0 $X=10096000 $Y=13552000
X5857 24 5615 ICV_19 $T=10112000 8448000 0 0 $X=10112000 $Y=8448000
X5858 24 5616 ICV_19 $T=10264000 5432000 0 0 $X=10264000 $Y=5432000
X5859 24 5617 ICV_19 $T=10392000 11696000 0 0 $X=10392000 $Y=11696000
X5860 24 5618 ICV_19 $T=10440000 4736000 0 0 $X=10440000 $Y=4736000
X5861 24 5619 ICV_19 $T=10480000 13088000 0 0 $X=10480000 $Y=13088000
X5862 24 5620 ICV_19 $T=10976000 6128000 0 0 $X=10976000 $Y=6128000
X5863 24 5621 ICV_19 $T=11024000 3808000 0 0 $X=11024000 $Y=3808000
X5864 24 5622 ICV_19 $T=11024000 4736000 0 0 $X=11024000 $Y=4736000
X5865 24 5623 ICV_19 $T=11128000 3576000 0 0 $X=11128000 $Y=3576000
X5866 24 5624 ICV_19 $T=11128000 7984000 0 0 $X=11128000 $Y=7984000
X5867 24 5625 ICV_19 $T=11240000 2416000 0 0 $X=11240000 $Y=2416000
X5868 24 4577 ICV_19 $T=11368000 1952000 0 0 $X=11368000 $Y=1952000
X5869 24 5626 ICV_19 $T=11472000 10304000 0 0 $X=11472000 $Y=10304000
X5870 24 5627 ICV_19 $T=11600000 9144000 0 0 $X=11600000 $Y=9144000
X5871 24 ICV_20 $T=584000 4272000 0 0 $X=584000 $Y=4272000
X5872 24 ICV_20 $T=688000 4040000 0 0 $X=688000 $Y=4040000
X5873 24 ICV_20 $T=944000 2880000 0 0 $X=944000 $Y=2880000
X5874 24 ICV_20 $T=1104000 96000 0 0 $X=1104000 $Y=96000
X5875 24 ICV_20 $T=1288000 792000 0 0 $X=1288000 $Y=792000
X5876 24 ICV_20 $T=3000000 560000 0 0 $X=3000000 $Y=560000
X5877 24 ICV_20 $T=3072000 328000 0 0 $X=3072000 $Y=328000
X5878 24 ICV_20 $T=11592000 7056000 0 0 $X=11592000 $Y=7056000
X5879 24 ICV_21 $T=4704000 1024000 1 180 $X=4520000 $Y=1024000
X5880 24 ICV_21 $T=6632000 6128000 1 180 $X=6448000 $Y=6128000
X5881 24 ICV_21 $T=8616000 2648000 1 180 $X=8432000 $Y=2648000
X5882 24 ICV_21 $T=9136000 2416000 1 180 $X=8952000 $Y=2416000
X5883 24 ICV_21 $T=9536000 6824000 1 180 $X=9352000 $Y=6824000
X5884 24 ICV_21 $T=10744000 10072000 1 180 $X=10560000 $Y=10072000
X5885 24 ICV_21 $T=11736000 7984000 1 180 $X=11552000 $Y=7984000
X5886 24 ICV_22 $T=559000 2184000 1 180 $X=496000 $Y=2184000
X5887 24 ICV_22 $T=791000 3808000 1 180 $X=728000 $Y=3808000
X5888 24 ICV_22 $T=1311000 2184000 1 180 $X=1248000 $Y=2184000
X5889 24 ICV_22 $T=1959000 1256000 1 180 $X=1896000 $Y=1256000
X5890 24 ICV_22 $T=2911000 560000 1 180 $X=2848000 $Y=560000
X5891 24 ICV_22 $T=11559000 6824000 1 180 $X=11496000 $Y=6824000
X5892 24 5628 ICV_23 $T=1312000 10536000 0 0 $X=1312000 $Y=10536000
X5893 24 5629 ICV_23 $T=1392000 10304000 0 0 $X=1392000 $Y=10304000
X5894 24 5630 ICV_23 $T=5408000 10536000 0 0 $X=5408000 $Y=10536000
X5895 24 5631 ICV_23 $T=5752000 10768000 0 0 $X=5752000 $Y=10768000
X5896 24 5329 ICV_23 $T=10960000 13552000 0 0 $X=10960000 $Y=13552000
X5897 24 5632 ICV_23 $T=11168000 12160000 0 0 $X=11168000 $Y=12160000
X5898 24 5633 ICV_23 $T=11448000 12160000 0 0 $X=11448000 $Y=12160000
X5899 24 ICV_24 $T=3160000 3576000 0 0 $X=3160000 $Y=3576000
X5900 24 ICV_24 $T=6152000 7520000 0 0 $X=6152000 $Y=7520000
X5901 24 ICV_24 $T=7024000 5896000 0 0 $X=7024000 $Y=5896000
X5902 24 ICV_24 $T=7680000 11000000 0 0 $X=7680000 $Y=11000000
X5903 24 ICV_24 $T=7880000 11928000 0 0 $X=7880000 $Y=11928000
X5904 24 ICV_24 $T=8608000 6592000 0 0 $X=8608000 $Y=6592000
X5905 24 ICV_24 $T=9168000 2416000 0 0 $X=9168000 $Y=2416000
X5906 24 ICV_24 $T=10424000 8448000 0 0 $X=10424000 $Y=8448000
X5907 24 ICV_24 $T=11448000 4504000 0 0 $X=11448000 $Y=4504000
X5908 24 ICV_25 $T=600000 1952000 0 0 $X=600000 $Y=1952000
X5909 24 ICV_25 $T=2032000 560000 0 0 $X=2032000 $Y=560000
X5910 24 ICV_25 $T=2696000 560000 0 0 $X=2696000 $Y=560000
X5911 24 ICV_25 $T=11424000 1720000 0 0 $X=11424000 $Y=1720000
X5912 24 oai32 $T=985000 3576000 1 180 $X=928000 $Y=3576000
X5913 24 oai32 $T=1001000 4040000 1 180 $X=944000 $Y=4040000
X5914 24 oai32 $T=1065000 4040000 1 180 $X=1008000 $Y=4040000
X5915 24 oai32 $T=1152000 3344000 0 0 $X=1152000 $Y=3344000
X5916 24 oai32 $T=1216000 3344000 0 0 $X=1216000 $Y=3344000
X5917 24 oai32 $T=1216000 3576000 0 0 $X=1216000 $Y=3576000
X5918 24 oai32 $T=1280000 3576000 0 0 $X=1280000 $Y=3576000
X5919 24 oai32 $T=1377000 4040000 1 180 $X=1320000 $Y=4040000
X5920 24 oai32 $T=1609000 4040000 1 180 $X=1552000 $Y=4040000
X5921 24 oai32 $T=2024000 3112000 0 0 $X=2024000 $Y=3112000
X5922 24 oai32 $T=10769000 1024000 1 180 $X=10712000 $Y=1024000
X5923 24 oai32 $T=10921000 1024000 1 180 $X=10864000 $Y=1024000
X5924 24 oai32 $T=10928000 1024000 0 0 $X=10928000 $Y=1024000
X5925 24 oai32 $T=11321000 6592000 1 180 $X=11264000 $Y=6592000
X5926 24 oai32 $T=11296000 1720000 0 0 $X=11296000 $Y=1720000
X5927 24 oai32 $T=11360000 6592000 0 0 $X=11360000 $Y=6592000
X5928 24 or04 $T=11393000 1488000 1 180 $X=11328000 $Y=1488000
X5929 24 5634 and02 $T=1529500 3112000 1 180 $X=1488000 $Y=3112000
X5930 24 5635 and02 $T=1568000 3112000 0 0 $X=1568000 $Y=3112000
X5931 24 5636 and02 $T=1793500 3112000 1 180 $X=1752000 $Y=3112000
X5932 24 5637 and02 $T=2440000 1952000 0 0 $X=2440000 $Y=1952000
X5933 24 5638 and02 $T=2456000 1720000 0 0 $X=2456000 $Y=1720000
X5934 24 5328 and02 $T=10712000 3112000 0 0 $X=10712000 $Y=3112000
X5935 24 5639 and02 $T=11288000 6824000 0 0 $X=11288000 $Y=6824000
X5936 24 ICV_26 $T=1288000 11928000 0 0 $X=1288000 $Y=11928000
X5937 24 ICV_26 $T=1808000 11232000 0 0 $X=1808000 $Y=11232000
X5938 24 ICV_26 $T=1920000 12624000 0 0 $X=1920000 $Y=12624000
X5939 24 ICV_26 $T=1960000 6592000 0 0 $X=1960000 $Y=6592000
X5940 24 ICV_26 $T=2200000 4968000 0 0 $X=2200000 $Y=4968000
X5941 24 ICV_26 $T=2240000 6592000 0 0 $X=2240000 $Y=6592000
X5942 24 ICV_26 $T=2328000 12624000 0 0 $X=2328000 $Y=12624000
X5943 24 ICV_26 $T=2936000 4272000 0 0 $X=2936000 $Y=4272000
X5944 24 ICV_26 $T=2952000 7288000 0 0 $X=2952000 $Y=7288000
X5945 24 ICV_26 $T=3208000 10072000 0 0 $X=3208000 $Y=10072000
X5946 24 ICV_26 $T=3352000 6824000 0 0 $X=3352000 $Y=6824000
X5947 24 ICV_26 $T=3800000 9376000 0 0 $X=3800000 $Y=9376000
X5948 24 ICV_26 $T=3936000 5432000 0 0 $X=3936000 $Y=5432000
X5949 24 ICV_26 $T=4200000 7520000 0 0 $X=4200000 $Y=7520000
X5950 24 ICV_26 $T=4232000 1720000 0 0 $X=4232000 $Y=1720000
X5951 24 ICV_26 $T=4504000 4040000 0 0 $X=4504000 $Y=4040000
X5952 24 ICV_26 $T=4536000 13088000 0 0 $X=4536000 $Y=13088000
X5953 24 ICV_26 $T=4560000 328000 0 0 $X=4560000 $Y=328000
X5954 24 ICV_26 $T=4712000 1256000 0 0 $X=4712000 $Y=1256000
X5955 24 ICV_26 $T=4760000 12160000 0 0 $X=4760000 $Y=12160000
X5956 24 ICV_26 $T=4832000 96000 0 0 $X=4832000 $Y=96000
X5957 24 ICV_26 $T=4832000 2416000 0 0 $X=4832000 $Y=2416000
X5958 24 ICV_26 $T=4880000 4272000 0 0 $X=4880000 $Y=4272000
X5959 24 ICV_26 $T=5008000 12160000 0 0 $X=5008000 $Y=12160000
X5960 24 ICV_26 $T=5256000 8448000 0 0 $X=5256000 $Y=8448000
X5961 24 ICV_26 $T=5304000 7056000 0 0 $X=5304000 $Y=7056000
X5962 24 ICV_26 $T=5344000 10072000 0 0 $X=5344000 $Y=10072000
X5963 24 ICV_26 $T=5368000 2880000 0 0 $X=5368000 $Y=2880000
X5964 24 ICV_26 $T=5664000 10304000 0 0 $X=5664000 $Y=10304000
X5965 24 ICV_26 $T=5688000 1720000 0 0 $X=5688000 $Y=1720000
X5966 24 ICV_26 $T=5744000 11928000 0 0 $X=5744000 $Y=11928000
X5967 24 ICV_26 $T=5808000 96000 0 0 $X=5808000 $Y=96000
X5968 24 ICV_26 $T=5808000 12392000 0 0 $X=5808000 $Y=12392000
X5969 24 ICV_26 $T=6104000 9144000 0 0 $X=6104000 $Y=9144000
X5970 24 ICV_26 $T=6112000 1488000 0 0 $X=6112000 $Y=1488000
X5971 24 ICV_26 $T=6128000 1024000 0 0 $X=6128000 $Y=1024000
X5972 24 ICV_26 $T=6152000 11928000 0 0 $X=6152000 $Y=11928000
X5973 24 ICV_26 $T=6152000 12160000 0 0 $X=6152000 $Y=12160000
X5974 24 ICV_26 $T=6168000 560000 0 0 $X=6168000 $Y=560000
X5975 24 ICV_26 $T=6168000 2416000 0 0 $X=6168000 $Y=2416000
X5976 24 ICV_26 $T=6192000 12624000 0 0 $X=6192000 $Y=12624000
X5977 24 ICV_26 $T=6416000 13320000 0 0 $X=6416000 $Y=13320000
X5978 24 ICV_26 $T=6432000 11928000 0 0 $X=6432000 $Y=11928000
X5979 24 ICV_26 $T=6504000 1952000 0 0 $X=6504000 $Y=1952000
X5980 24 ICV_26 $T=6672000 4272000 0 0 $X=6672000 $Y=4272000
X5981 24 ICV_26 $T=6696000 5432000 0 0 $X=6696000 $Y=5432000
X5982 24 ICV_26 $T=6808000 3344000 0 0 $X=6808000 $Y=3344000
X5983 24 ICV_26 $T=7112000 2416000 0 0 $X=7112000 $Y=2416000
X5984 24 ICV_26 $T=7656000 9840000 0 0 $X=7656000 $Y=9840000
X5985 24 ICV_26 $T=7664000 4272000 0 0 $X=7664000 $Y=4272000
X5986 24 ICV_26 $T=7744000 8680000 0 0 $X=7744000 $Y=8680000
X5987 24 ICV_26 $T=7768000 8912000 0 0 $X=7768000 $Y=8912000
X5988 24 ICV_26 $T=7776000 3576000 0 0 $X=7776000 $Y=3576000
X5989 24 ICV_26 $T=7808000 4040000 0 0 $X=7808000 $Y=4040000
X5990 24 ICV_26 $T=8320000 11696000 0 0 $X=8320000 $Y=11696000
X5991 24 ICV_26 $T=8488000 96000 0 0 $X=8488000 $Y=96000
X5992 24 ICV_26 $T=8536000 8448000 0 0 $X=8536000 $Y=8448000
X5993 24 ICV_26 $T=9080000 2880000 0 0 $X=9080000 $Y=2880000
X5994 24 ICV_26 $T=9112000 1256000 0 0 $X=9112000 $Y=1256000
X5995 24 ICV_26 $T=9728000 3112000 0 0 $X=9728000 $Y=3112000
X5996 24 ICV_26 $T=10240000 3344000 0 0 $X=10240000 $Y=3344000
X5997 24 ICV_26 $T=10504000 6824000 0 0 $X=10504000 $Y=6824000
X5998 24 ICV_26 $T=10888000 12624000 0 0 $X=10888000 $Y=12624000
X5999 24 ICV_26 $T=11064000 5664000 0 0 $X=11064000 $Y=5664000
X6000 24 ICV_26 $T=11112000 4040000 0 0 $X=11112000 $Y=4040000
X6001 24 nor02_2x $T=448000 8448000 0 0 $X=448000 $Y=8448000
X6002 24 nor02_2x $T=688000 8912000 0 0 $X=688000 $Y=8912000
X6003 24 nor02_2x $T=696000 8680000 0 0 $X=696000 $Y=8680000
X6004 24 nor02_2x $T=1473000 9840000 1 180 $X=1440000 $Y=9840000
X6005 24 nor02_2x $T=1616000 9840000 0 0 $X=1616000 $Y=9840000
X6006 24 nor02_2x $T=1752000 2184000 0 0 $X=1752000 $Y=2184000
X6007 24 nor02_2x $T=1776000 10072000 0 0 $X=1776000 $Y=10072000
X6008 24 nor02_2x $T=2129000 1720000 1 180 $X=2096000 $Y=1720000
X6009 24 nor02_2x $T=2344000 1952000 0 0 $X=2344000 $Y=1952000
X6010 24 nor02_2x $T=2848000 2648000 0 0 $X=2848000 $Y=2648000
X6011 24 nor02_2x $T=10528000 1256000 0 0 $X=10528000 $Y=1256000
X6012 24 nor02_2x $T=11081000 1488000 1 180 $X=11048000 $Y=1488000
X6013 24 ICV_27 $T=152000 10536000 0 0 $X=152000 $Y=10536000
X6014 24 ICV_27 $T=152000 11696000 0 0 $X=152000 $Y=11696000
X6015 24 ICV_27 $T=216000 11232000 0 0 $X=216000 $Y=11232000
X6016 24 ICV_27 $T=432000 13552000 0 0 $X=432000 $Y=13552000
X6017 24 ICV_27 $T=1104000 12160000 0 0 $X=1104000 $Y=12160000
X6018 24 ICV_27 $T=1360000 11464000 0 0 $X=1360000 $Y=11464000
X6019 24 ICV_27 $T=1392000 13320000 0 0 $X=1392000 $Y=13320000
X6020 24 ICV_27 $T=1416000 12856000 0 0 $X=1416000 $Y=12856000
X6021 24 ICV_27 $T=2224000 8216000 0 0 $X=2224000 $Y=8216000
X6022 24 ICV_27 $T=2384000 5896000 0 0 $X=2384000 $Y=5896000
X6023 24 ICV_27 $T=2688000 5432000 0 0 $X=2688000 $Y=5432000
X6024 24 ICV_27 $T=2992000 6128000 0 0 $X=2992000 $Y=6128000
X6025 24 ICV_27 $T=3184000 5432000 0 0 $X=3184000 $Y=5432000
X6026 24 ICV_27 $T=3192000 2648000 0 0 $X=3192000 $Y=2648000
X6027 24 ICV_27 $T=3280000 4272000 0 0 $X=3280000 $Y=4272000
X6028 24 ICV_27 $T=3312000 3112000 0 0 $X=3312000 $Y=3112000
X6029 24 ICV_27 $T=3496000 12856000 0 0 $X=3496000 $Y=12856000
X6030 24 ICV_27 $T=3752000 1488000 0 0 $X=3752000 $Y=1488000
X6031 24 ICV_27 $T=3784000 8912000 0 0 $X=3784000 $Y=8912000
X6032 24 ICV_27 $T=3936000 8680000 0 0 $X=3936000 $Y=8680000
X6033 24 ICV_27 $T=3976000 4736000 0 0 $X=3976000 $Y=4736000
X6034 24 ICV_27 $T=4680000 3344000 0 0 $X=4680000 $Y=3344000
X6035 24 ICV_27 $T=4744000 3576000 0 0 $X=4744000 $Y=3576000
X6036 24 ICV_27 $T=4760000 11464000 0 0 $X=4760000 $Y=11464000
X6037 24 ICV_27 $T=5432000 2648000 0 0 $X=5432000 $Y=2648000
X6038 24 ICV_27 $T=5528000 4040000 0 0 $X=5528000 $Y=4040000
X6039 24 ICV_27 $T=5544000 3576000 0 0 $X=5544000 $Y=3576000
X6040 24 ICV_27 $T=7048000 8912000 0 0 $X=7048000 $Y=8912000
X6041 24 ICV_27 $T=7144000 2648000 0 0 $X=7144000 $Y=2648000
X6042 24 ICV_27 $T=7264000 10304000 0 0 $X=7264000 $Y=10304000
X6043 24 ICV_27 $T=7576000 7752000 0 0 $X=7576000 $Y=7752000
X6044 24 ICV_27 $T=7664000 9376000 0 0 $X=7664000 $Y=9376000
X6045 24 ICV_27 $T=7728000 3808000 0 0 $X=7728000 $Y=3808000
X6046 24 ICV_27 $T=8360000 3576000 0 0 $X=8360000 $Y=3576000
X6047 24 ICV_27 $T=8560000 1256000 0 0 $X=8560000 $Y=1256000
X6048 24 ICV_27 $T=8632000 4504000 0 0 $X=8632000 $Y=4504000
X6049 24 ICV_27 $T=8848000 7520000 0 0 $X=8848000 $Y=7520000
X6050 24 ICV_27 $T=9248000 10304000 0 0 $X=9248000 $Y=10304000
X6051 24 ICV_27 $T=9272000 10536000 0 0 $X=9272000 $Y=10536000
X6052 24 ICV_27 $T=9320000 10768000 0 0 $X=9320000 $Y=10768000
X6053 24 ICV_27 $T=9368000 11696000 0 0 $X=9368000 $Y=11696000
X6054 24 ICV_27 $T=9392000 9840000 0 0 $X=9392000 $Y=9840000
X6055 24 ICV_27 $T=9704000 7288000 0 0 $X=9704000 $Y=7288000
X6056 24 ICV_27 $T=10856000 9608000 0 0 $X=10856000 $Y=9608000
X6057 24 ICV_27 $T=10904000 4968000 0 0 $X=10904000 $Y=4968000
X6058 24 ICV_27 $T=10952000 4504000 0 0 $X=10952000 $Y=4504000
X6059 24 ICV_28 $T=336000 7288000 1 180 $X=152000 $Y=7288000
X6060 24 ICV_28 $T=3208000 7984000 1 180 $X=3024000 $Y=7984000
X6061 24 ICV_28 $T=4008000 11464000 1 180 $X=3824000 $Y=11464000
X6062 24 ICV_28 $T=7176000 2184000 1 180 $X=6992000 $Y=2184000
X6063 24 ICV_28 $T=7808000 13088000 1 180 $X=7624000 $Y=13088000
X6064 24 ICV_28 $T=8768000 1720000 1 180 $X=8584000 $Y=1720000
X6065 24 ICV_28 $T=11096000 5896000 1 180 $X=10912000 $Y=5896000
X6066 24 ao22 $T=10864000 560000 0 0 $X=10864000 $Y=560000
X6067 24 ICV_29 $T=1440000 13088000 0 0 $X=1440000 $Y=13088000
X6068 24 ICV_29 $T=2200000 7288000 0 0 $X=2200000 $Y=7288000
X6069 24 ICV_29 $T=3304000 4504000 0 0 $X=3304000 $Y=4504000
X6070 24 ICV_29 $T=3592000 3576000 0 0 $X=3592000 $Y=3576000
X6071 24 ICV_29 $T=3744000 11000000 0 0 $X=3744000 $Y=11000000
X6072 24 ICV_29 $T=6888000 2880000 0 0 $X=6888000 $Y=2880000
X6073 24 ICV_29 $T=9368000 6128000 0 0 $X=9368000 $Y=6128000
X6074 24 ICV_29 $T=10432000 10304000 0 0 $X=10432000 $Y=10304000
X6075 24 ICV_29 $T=10824000 6360000 0 0 $X=10824000 $Y=6360000
X6076 24 aoi221 $T=10881500 1488000 1 180 $X=10816000 $Y=1488000
X6077 24 5640 oai21 $T=897000 11928000 1 180 $X=856000 $Y=11928000
X6078 24 5641 oai21 $T=904000 11928000 0 0 $X=904000 $Y=11928000
X6079 24 5642 oai21 $T=1049000 11928000 1 180 $X=1008000 $Y=11928000
X6080 24 5643 oai21 $T=1145000 2648000 1 180 $X=1104000 $Y=2648000
X6081 24 5644 oai21 $T=1193000 3112000 1 180 $X=1152000 $Y=3112000
X6082 24 5645 oai21 $T=1200000 3112000 0 0 $X=1200000 $Y=3112000
X6083 24 5646 oai21 $T=1328000 3112000 0 0 $X=1328000 $Y=3112000
X6084 24 5647 oai21 $T=1472000 7520000 0 0 $X=1472000 $Y=7520000
X6085 24 5648 oai21 $T=1520000 7520000 0 0 $X=1520000 $Y=7520000
X6086 24 5649 oai21 $T=1536000 6128000 0 0 $X=1536000 $Y=6128000
X6087 24 5650 oai21 $T=1560000 7752000 0 0 $X=1560000 $Y=7752000
X6088 24 5651 oai21 $T=1584000 6128000 0 0 $X=1584000 $Y=6128000
X6089 24 5652 oai21 $T=1608000 5432000 0 0 $X=1608000 $Y=5432000
X6090 24 5653 oai21 $T=1632000 11000000 0 0 $X=1632000 $Y=11000000
X6091 24 5654 oai21 $T=1640000 7520000 0 0 $X=1640000 $Y=7520000
X6092 24 5655 oai21 $T=1656000 5432000 0 0 $X=1656000 $Y=5432000
X6093 24 5656 oai21 $T=1968000 2880000 0 0 $X=1968000 $Y=2880000
X6094 24 5657 oai21 $T=2369000 3112000 1 180 $X=2328000 $Y=3112000
X6095 24 5658 oai21 $T=2409000 2880000 1 180 $X=2368000 $Y=2880000
X6096 24 5659 oai21 $T=2488000 3112000 0 0 $X=2488000 $Y=3112000
X6097 24 5660 oai21 $T=2561000 4272000 1 180 $X=2520000 $Y=4272000
X6098 24 5661 oai21 $T=2569000 4504000 1 180 $X=2528000 $Y=4504000
X6099 24 5662 oai21 $T=2560000 2880000 0 0 $X=2560000 $Y=2880000
X6100 24 5663 oai21 $T=2576000 4736000 0 0 $X=2576000 $Y=4736000
X6101 24 5664 oai21 $T=2608000 2880000 0 0 $X=2608000 $Y=2880000
X6102 24 5665 oai21 $T=2888000 2648000 0 0 $X=2888000 $Y=2648000
X6103 24 5666 oai21 $T=3313000 9144000 1 180 $X=3272000 $Y=9144000
X6104 24 5667 oai21 $T=3425000 12160000 1 180 $X=3384000 $Y=12160000
X6105 24 5668 oai21 $T=3433000 12392000 1 180 $X=3392000 $Y=12392000
X6106 24 5669 oai21 $T=3665000 12160000 1 180 $X=3624000 $Y=12160000
X6107 24 5670 oai21 $T=3728000 5200000 0 0 $X=3728000 $Y=5200000
X6108 24 5671 oai21 $T=3769000 12160000 1 180 $X=3728000 $Y=12160000
X6109 24 5672 oai21 $T=3785000 12392000 1 180 $X=3744000 $Y=12392000
X6110 24 5673 oai21 $T=3817000 5200000 1 180 $X=3776000 $Y=5200000
X6111 24 5674 oai21 $T=3865000 5200000 1 180 $X=3824000 $Y=5200000
X6112 24 5675 oai21 $T=3889000 12392000 1 180 $X=3848000 $Y=12392000
X6113 24 5676 oai21 $T=3913000 7752000 1 180 $X=3872000 $Y=7752000
X6114 24 5677 oai21 $T=3921000 9608000 1 180 $X=3880000 $Y=9608000
X6115 24 5678 oai21 $T=3937000 12392000 1 180 $X=3896000 $Y=12392000
X6116 24 5679 oai21 $T=3969000 9608000 1 180 $X=3928000 $Y=9608000
X6117 24 5680 oai21 $T=3985000 9144000 1 180 $X=3944000 $Y=9144000
X6118 24 5681 oai21 $T=3993000 9840000 1 180 $X=3952000 $Y=9840000
X6119 24 5682 oai21 $T=4105000 12160000 1 180 $X=4064000 $Y=12160000
X6120 24 5683 oai21 $T=4280000 9608000 0 0 $X=4280000 $Y=9608000
X6121 24 5684 oai21 $T=4336000 4272000 0 0 $X=4336000 $Y=4272000
X6122 24 5685 oai21 $T=4409000 11000000 1 180 $X=4368000 $Y=11000000
X6123 24 5686 oai21 $T=4600000 792000 0 0 $X=4600000 $Y=792000
X6124 24 5687 oai21 $T=4648000 792000 0 0 $X=4648000 $Y=792000
X6125 24 5688 oai21 $T=4689000 7752000 1 180 $X=4648000 $Y=7752000
X6126 24 5325 oai21 $T=4664000 1256000 0 0 $X=4664000 $Y=1256000
X6127 24 5689 oai21 $T=4664000 2184000 0 0 $X=4664000 $Y=2184000
X6128 24 5690 oai21 $T=4688000 1952000 0 0 $X=4688000 $Y=1952000
X6129 24 5691 oai21 $T=4761000 7520000 1 180 $X=4720000 $Y=7520000
X6130 24 5692 oai21 $T=4752000 792000 0 0 $X=4752000 $Y=792000
X6131 24 5693 oai21 $T=4768000 2184000 0 0 $X=4768000 $Y=2184000
X6132 24 5694 oai21 $T=5065000 10768000 1 180 $X=5024000 $Y=10768000
X6133 24 5695 oai21 $T=5089000 6360000 1 180 $X=5048000 $Y=6360000
X6134 24 5696 oai21 $T=5072000 8912000 0 0 $X=5072000 $Y=8912000
X6135 24 5697 oai21 $T=5225000 11232000 1 180 $X=5184000 $Y=11232000
X6136 24 5698 oai21 $T=5361000 5664000 1 180 $X=5320000 $Y=5664000
X6137 24 5699 oai21 $T=5473000 6592000 1 180 $X=5432000 $Y=6592000
X6138 24 5700 oai21 $T=5569000 4736000 1 180 $X=5528000 $Y=4736000
X6139 24 5701 oai21 $T=6208000 3808000 0 0 $X=6208000 $Y=3808000
X6140 24 5702 oai21 $T=6569000 5200000 1 180 $X=6528000 $Y=5200000
X6141 24 5703 oai21 $T=6625000 3576000 1 180 $X=6584000 $Y=3576000
X6142 24 5704 oai21 $T=6776000 12160000 0 0 $X=6776000 $Y=12160000
X6143 24 5705 oai21 $T=6880000 1024000 0 0 $X=6880000 $Y=1024000
X6144 24 4099 oai21 $T=6904000 10304000 0 0 $X=6904000 $Y=10304000
X6145 24 5706 oai21 $T=6944000 8912000 0 0 $X=6944000 $Y=8912000
X6146 24 5707 oai21 $T=6993000 4504000 1 180 $X=6952000 $Y=4504000
X6147 24 5708 oai21 $T=7065000 12160000 1 180 $X=7024000 $Y=12160000
X6148 24 5709 oai21 $T=7097000 4504000 1 180 $X=7056000 $Y=4504000
X6149 24 5710 oai21 $T=7153000 7288000 1 180 $X=7112000 $Y=7288000
X6150 24 5711 oai21 $T=7177000 12160000 1 180 $X=7136000 $Y=12160000
X6151 24 5712 oai21 $T=7216000 12160000 0 0 $X=7216000 $Y=12160000
X6152 24 5327 oai21 $T=7280000 7056000 0 0 $X=7280000 $Y=7056000
X6153 24 5713 oai21 $T=7288000 1024000 0 0 $X=7288000 $Y=1024000
X6154 24 5714 oai21 $T=7377000 4504000 1 180 $X=7336000 $Y=4504000
X6155 24 5715 oai21 $T=7424000 1024000 0 0 $X=7424000 $Y=1024000
X6156 24 5716 oai21 $T=7696000 5896000 0 0 $X=7696000 $Y=5896000
X6157 24 5717 oai21 $T=7760000 11696000 0 0 $X=7760000 $Y=11696000
X6158 24 5718 oai21 $T=7776000 5432000 0 0 $X=7776000 $Y=5432000
X6159 24 5719 oai21 $T=7920000 2880000 0 0 $X=7920000 $Y=2880000
X6160 24 5720 oai21 $T=8032000 2880000 0 0 $X=8032000 $Y=2880000
X6161 24 5721 oai21 $T=8048000 1720000 0 0 $X=8048000 $Y=1720000
X6162 24 5722 oai21 $T=8152000 5200000 0 0 $X=8152000 $Y=5200000
X6163 24 5723 oai21 $T=8248000 2880000 0 0 $X=8248000 $Y=2880000
X6164 24 5724 oai21 $T=8264000 560000 0 0 $X=8264000 $Y=560000
X6165 24 5725 oai21 $T=8280000 1952000 0 0 $X=8280000 $Y=1952000
X6166 24 5726 oai21 $T=8304000 8680000 0 0 $X=8304000 $Y=8680000
X6167 24 5727 oai21 $T=8336000 4968000 0 0 $X=8336000 $Y=4968000
X6168 24 5728 oai21 $T=8416000 792000 0 0 $X=8416000 $Y=792000
X6169 24 2344 oai21 $T=8736000 4736000 0 0 $X=8736000 $Y=4736000
X6170 24 5729 oai21 $T=8929000 12624000 1 180 $X=8888000 $Y=12624000
X6171 24 5730 oai21 $T=8936000 1024000 0 0 $X=8936000 $Y=1024000
X6172 24 5731 oai21 $T=8977000 12624000 1 180 $X=8936000 $Y=12624000
X6173 24 5732 oai21 $T=8968000 11928000 0 0 $X=8968000 $Y=11928000
X6174 24 2346 oai21 $T=9152000 3808000 0 0 $X=9152000 $Y=3808000
X6175 24 5733 oai21 $T=9417000 7288000 1 180 $X=9376000 $Y=7288000
X6176 24 5734 oai21 $T=9416000 9376000 0 0 $X=9416000 $Y=9376000
X6177 24 5735 oai21 $T=9432000 12392000 0 0 $X=9432000 $Y=12392000
X6178 24 5736 oai21 $T=10072000 10304000 0 0 $X=10072000 $Y=10304000
X6179 24 5737 oai21 $T=10104000 9376000 0 0 $X=10104000 $Y=9376000
X6180 24 5738 oai21 $T=10312000 4504000 0 0 $X=10312000 $Y=4504000
X6181 24 5739 oai21 $T=10392000 11000000 0 0 $X=10392000 $Y=11000000
X6182 24 5740 oai21 $T=10416000 3808000 0 0 $X=10416000 $Y=3808000
X6183 24 5741 oai21 $T=10465000 8680000 1 180 $X=10424000 $Y=8680000
X6184 24 5742 oai21 $T=10440000 11000000 0 0 $X=10440000 $Y=11000000
X6185 24 5743 oai21 $T=10480000 3576000 0 0 $X=10480000 $Y=3576000
X6186 24 5744 oai21 $T=10512000 9376000 0 0 $X=10512000 $Y=9376000
X6187 24 5745 oai21 $T=10617000 3808000 1 180 $X=10576000 $Y=3808000
X6188 24 5746 oai21 $T=10600000 4040000 0 0 $X=10600000 $Y=4040000
X6189 24 5747 oai21 $T=10632000 7984000 0 0 $X=10632000 $Y=7984000
X6190 24 5748 oai21 $T=10705000 6360000 1 180 $X=10664000 $Y=6360000
X6191 24 5749 oai21 $T=10688000 9608000 0 0 $X=10688000 $Y=9608000
X6192 24 5750 oai21 $T=10704000 5896000 0 0 $X=10704000 $Y=5896000
X6193 24 5751 oai21 $T=10712000 4272000 0 0 $X=10712000 $Y=4272000
X6194 24 5752 oai21 $T=10712000 7984000 0 0 $X=10712000 $Y=7984000
X6195 24 5753 oai21 $T=10793000 10768000 1 180 $X=10752000 $Y=10768000
X6196 24 5754 oai21 $T=10760000 4272000 0 0 $X=10760000 $Y=4272000
X6197 24 4101 oai21 $T=10760000 7752000 0 0 $X=10760000 $Y=7752000
X6198 24 5755 oai21 $T=10776000 6360000 0 0 $X=10776000 $Y=6360000
X6199 24 5756 oai21 $T=10784000 11000000 0 0 $X=10784000 $Y=11000000
X6200 24 5757 oai21 $T=10808000 5896000 0 0 $X=10808000 $Y=5896000
X6201 24 nor03_2x $T=289000 3112000 1 180 $X=248000 $Y=3112000
X6202 24 nor03_2x $T=337000 3112000 1 180 $X=296000 $Y=3112000
X6203 24 nor03_2x $T=1344000 3344000 0 0 $X=1344000 $Y=3344000
X6204 24 nor03_2x $T=1441000 2648000 1 180 $X=1400000 $Y=2648000
X6205 24 nor03_2x $T=1496000 2648000 0 0 $X=1496000 $Y=2648000
X6206 24 nor03_2x $T=1665000 2880000 1 180 $X=1624000 $Y=2880000
X6207 24 nor03_2x $T=1680000 2416000 0 0 $X=1680000 $Y=2416000
X6208 24 nor03_2x $T=1801000 2880000 1 180 $X=1760000 $Y=2880000
X6209 24 nor03_2x $T=1825000 2648000 1 180 $X=1784000 $Y=2648000
X6210 24 nor03_2x $T=1888000 2648000 0 0 $X=1888000 $Y=2648000
X6211 24 nor03_2x $T=2032000 2416000 0 0 $X=2032000 $Y=2416000
X6212 24 nor03_2x $T=2121000 2416000 1 180 $X=2080000 $Y=2416000
X6213 24 nor03_2x $T=2225000 2648000 1 180 $X=2184000 $Y=2648000
X6214 24 nor03_2x $T=2345000 2184000 1 180 $X=2304000 $Y=2184000
X6215 24 nor03_2x $T=2464000 2184000 0 0 $X=2464000 $Y=2184000
X6216 24 nor03_2x $T=10377000 1488000 1 180 $X=10336000 $Y=1488000
X6217 24 nor03_2x $T=10585000 1488000 1 180 $X=10544000 $Y=1488000
X6218 24 nor03_2x $T=10808000 1256000 0 0 $X=10808000 $Y=1256000
X6219 24 inv04 $T=328000 4272000 0 0 $X=328000 $Y=4272000
X6220 24 inv04 $T=537000 3576000 1 180 $X=504000 $Y=3576000
X6221 24 inv04 $T=1601000 11696000 1 180 $X=1568000 $Y=11696000
X6222 24 inv04 $T=10776000 1488000 0 0 $X=10776000 $Y=1488000
X6223 24 aoi21 $T=193000 3112000 1 180 $X=152000 $Y=3112000
X6224 24 aoi21 $T=200000 3112000 0 0 $X=200000 $Y=3112000
X6225 24 aoi21 $T=1056000 3112000 0 0 $X=1056000 $Y=3112000
X6226 24 aoi21 $T=1104000 3112000 0 0 $X=1104000 $Y=3112000
X6227 24 aoi21 $T=1321000 3112000 1 180 $X=1280000 $Y=3112000
X6228 24 aoi21 $T=1440000 3344000 0 0 $X=1440000 $Y=3344000
X6229 24 aoi21 $T=1448000 2648000 0 0 $X=1448000 $Y=2648000
X6230 24 aoi21 $T=1456000 4040000 0 0 $X=1456000 $Y=4040000
X6231 24 aoi21 $T=1504000 4040000 0 0 $X=1504000 $Y=4040000
X6232 24 aoi21 $T=1536000 3344000 0 0 $X=1536000 $Y=3344000
X6233 24 aoi21 $T=1576000 2648000 0 0 $X=1576000 $Y=2648000
X6234 24 aoi21 $T=1617000 2880000 1 180 $X=1576000 $Y=2880000
X6235 24 aoi21 $T=2296000 1952000 0 0 $X=2296000 $Y=1952000
X6236 24 aoi21 $T=2384000 2184000 0 0 $X=2384000 $Y=2184000
X6237 24 aoi21 $T=2408000 1720000 0 0 $X=2408000 $Y=1720000
X6238 24 aoi21 $T=2512000 2184000 0 0 $X=2512000 $Y=2184000
X6239 24 aoi21 $T=2737000 2880000 1 180 $X=2696000 $Y=2880000
X6240 24 aoi21 $T=10769000 1256000 1 180 $X=10728000 $Y=1256000
X6241 24 ICV_30 $T=1880000 4504000 0 0 $X=1880000 $Y=4504000
X6242 24 ICV_30 $T=4104000 4272000 0 0 $X=4104000 $Y=4272000
X6243 24 ICV_30 $T=4520000 2648000 0 0 $X=4520000 $Y=2648000
X6244 24 ICV_30 $T=6664000 8216000 0 0 $X=6664000 $Y=8216000
X6245 24 ICV_30 $T=7056000 10768000 0 0 $X=7056000 $Y=10768000
X6246 24 ICV_30 $T=7064000 7984000 0 0 $X=7064000 $Y=7984000
X6247 24 ICV_30 $T=7816000 1720000 0 0 $X=7816000 $Y=1720000
X6248 24 ICV_30 $T=9168000 1952000 0 0 $X=9168000 $Y=1952000
X6249 24 ICV_30 $T=10552000 11000000 0 0 $X=10552000 $Y=11000000
X6250 24 ICV_31 $T=496000 7752000 0 0 $X=496000 $Y=7752000
X6251 24 ICV_31 $T=2472000 13320000 0 0 $X=2472000 $Y=13320000
X6252 24 ICV_31 $T=3152000 12392000 0 0 $X=3152000 $Y=12392000
X6253 24 ICV_31 $T=4056000 792000 0 0 $X=4056000 $Y=792000
X6254 24 ICV_31 $T=4152000 3808000 0 0 $X=4152000 $Y=3808000
X6255 24 ICV_31 $T=4832000 8680000 0 0 $X=4832000 $Y=8680000
X6256 24 ICV_31 $T=5288000 4736000 0 0 $X=5288000 $Y=4736000
X6257 24 ICV_31 $T=5752000 7752000 0 0 $X=5752000 $Y=7752000
X6258 24 ICV_31 $T=6608000 11464000 0 0 $X=6608000 $Y=11464000
X6259 24 ICV_31 $T=6864000 3576000 0 0 $X=6864000 $Y=3576000
X6260 24 ICV_31 $T=7632000 5200000 0 0 $X=7632000 $Y=5200000
X6261 24 ICV_31 $T=10128000 2648000 0 0 $X=10128000 $Y=2648000
X6262 24 ICV_31 $T=10280000 11232000 0 0 $X=10280000 $Y=11232000
X6263 24 ICV_31 $T=10448000 9608000 0 0 $X=10448000 $Y=9608000
X6264 24 ICV_32 $T=3680000 1720000 0 0 $X=3680000 $Y=1720000
X6265 24 ICV_32 $T=6600000 1256000 0 0 $X=6600000 $Y=1256000
X6266 24 ICV_32 $T=7408000 11464000 0 0 $X=7408000 $Y=11464000
X6267 24 ICV_32 $T=7448000 10536000 0 0 $X=7448000 $Y=10536000
X6268 24 ICV_32 $T=10056000 1720000 0 0 $X=10056000 $Y=1720000
X6269 24 ICV_33 $T=3552000 8912000 0 0 $X=3552000 $Y=8912000
X6270 24 ICV_33 $T=4448000 7288000 0 0 $X=4448000 $Y=7288000
X6271 24 ICV_33 $T=4816000 8216000 0 0 $X=4816000 $Y=8216000
X6272 24 ICV_33 $T=6544000 2648000 0 0 $X=6544000 $Y=2648000
X6273 24 ICV_33 $T=9184000 9376000 0 0 $X=9184000 $Y=9376000
X6274 24 ICV_33 $T=9936000 5432000 0 0 $X=9936000 $Y=5432000
X6275 24 5758 ICV_34 $T=2992000 4040000 0 0 $X=2992000 $Y=4040000
X6276 24 5759 ICV_34 $T=5104000 13552000 0 0 $X=5104000 $Y=13552000
X6277 24 5760 ICV_34 $T=6832000 7752000 0 0 $X=6832000 $Y=7752000
X6278 24 2343 ICV_34 $T=7728000 3344000 0 0 $X=7728000 $Y=3344000
X6279 24 5761 ICV_34 $T=9064000 11000000 0 0 $X=9064000 $Y=11000000
X6280 24 5762 ICV_34 $T=9120000 7752000 0 0 $X=9120000 $Y=7752000
X6281 24 5763 nor04 $T=1017000 3808000 1 180 $X=968000 $Y=3808000
X6282 24 5764 nor04 $T=2384000 1952000 0 0 $X=2384000 $Y=1952000
X6283 24 5765 nor04 $T=3568000 12160000 0 0 $X=3568000 $Y=12160000
X6284 24 2315 nor04 $T=3704000 7984000 0 0 $X=3704000 $Y=7984000
X6285 24 2319 nor04 $T=4696000 1720000 0 0 $X=4696000 $Y=1720000
X6286 24 2321 nor04 $T=4768000 6592000 0 0 $X=4768000 $Y=6592000
X6287 24 2329 nor04 $T=6328000 792000 0 0 $X=6328000 $Y=792000
X6288 24 5766 nor04 $T=7088000 8680000 0 0 $X=7088000 $Y=8680000
X6289 24 5767 nor04 $T=7104000 4504000 0 0 $X=7104000 $Y=4504000
X6290 24 5768 nor04 $T=7777000 4968000 1 180 $X=7728000 $Y=4968000
X6291 24 ICV_35 $T=2416000 8680000 1 180 $X=2232000 $Y=8680000
X6292 24 ICV_35 $T=4648000 6360000 1 180 $X=4464000 $Y=6360000
X6293 24 ICV_35 $T=4848000 10072000 1 180 $X=4664000 $Y=10072000
X6294 24 ICV_35 $T=5864000 6128000 1 180 $X=5680000 $Y=6128000
X6295 24 ICV_35 $T=6008000 1952000 1 180 $X=5824000 $Y=1952000
X6296 24 ICV_35 $T=6304000 7984000 1 180 $X=6120000 $Y=7984000
X6297 24 ICV_35 $T=7192000 6360000 1 180 $X=7008000 $Y=6360000
X6298 24 ICV_35 $T=7760000 3112000 1 180 $X=7576000 $Y=3112000
X6299 5769 24 or02 $T=2144000 1952000 0 0 $X=2144000 $Y=1952000
X6300 2325 24 or02 $T=5696000 96000 0 0 $X=5696000 $Y=96000
X6301 24 5770 or03 $T=1720000 11928000 0 0 $X=1720000 $Y=11928000
X6302 24 5771 or03 $T=1728000 11696000 0 0 $X=1728000 $Y=11696000
X6303 24 5772 or03 $T=1824000 11696000 0 0 $X=1824000 $Y=11696000
X6304 24 5773 or03 $T=1880000 11696000 0 0 $X=1880000 $Y=11696000
X6305 24 5774 or03 $T=1896000 11928000 0 0 $X=1896000 $Y=11928000
X6306 24 5775 or03 $T=1987000 2648000 1 180 $X=1936000 $Y=2648000
X6307 24 5776 or03 $T=1936000 11696000 0 0 $X=1936000 $Y=11696000
X6308 24 5777 or03 $T=1952000 11928000 0 0 $X=1952000 $Y=11928000
X6309 24 5778 or03 $T=2043000 11696000 1 180 $X=1992000 $Y=11696000
X6310 24 5779 or03 $T=2088000 11696000 0 0 $X=2088000 $Y=11696000
X6311 24 5780 or03 $T=2096000 11464000 0 0 $X=2096000 $Y=11464000
X6312 24 5781 or03 $T=2152000 11464000 0 0 $X=2152000 $Y=11464000
X6313 24 5782 or03 $T=2227000 11696000 1 180 $X=2176000 $Y=11696000
X6314 24 5783 or03 $T=2208000 11464000 0 0 $X=2208000 $Y=11464000
X6315 24 5784 or03 $T=2264000 11464000 0 0 $X=2264000 $Y=11464000
X6316 24 5785 or03 $T=2320000 11464000 0 0 $X=2320000 $Y=11464000
X6317 24 5786 or03 $T=2376000 11464000 0 0 $X=2376000 $Y=11464000
X6318 24 5787 or03 $T=2416000 2880000 0 0 $X=2416000 $Y=2880000
X6319 24 5788 or03 $T=2432000 11928000 0 0 $X=2432000 $Y=11928000
X6320 24 5789 or03 $T=2488000 11928000 0 0 $X=2488000 $Y=11928000
X6321 24 5790 or03 $T=2555000 2880000 1 180 $X=2504000 $Y=2880000
X6322 24 5791 or03 $T=2544000 11696000 0 0 $X=2544000 $Y=11696000
X6323 24 5792 or03 $T=2635000 11928000 1 180 $X=2584000 $Y=11928000
X6324 24 5793 or03 $T=2683000 11696000 1 180 $X=2632000 $Y=11696000
X6325 24 5794 or03 $T=2691000 11928000 1 180 $X=2640000 $Y=11928000
X6326 24 5795 or03 $T=2696000 11928000 0 0 $X=2696000 $Y=11928000
X6327 24 5796 or03 $T=2720000 11696000 0 0 $X=2720000 $Y=11696000
X6328 24 5797 or03 $T=2800000 11928000 0 0 $X=2800000 $Y=11928000
X6329 24 5798 or03 $T=2867000 11464000 1 180 $X=2816000 $Y=11464000
X6330 24 5799 or03 $T=2867000 11696000 1 180 $X=2816000 $Y=11696000
X6331 24 5800 or03 $T=2875000 11000000 1 180 $X=2824000 $Y=11000000
X6332 24 5801 or03 $T=2875000 11232000 1 180 $X=2824000 $Y=11232000
X6333 24 5802 or03 $T=2907000 11928000 1 180 $X=2856000 $Y=11928000
X6334 24 5803 or03 $T=2923000 11696000 1 180 $X=2872000 $Y=11696000
X6335 24 5804 or03 $T=2931000 11000000 1 180 $X=2880000 $Y=11000000
X6336 24 5805 or03 $T=2880000 11232000 0 0 $X=2880000 $Y=11232000
X6337 24 5806 or03 $T=2963000 11928000 1 180 $X=2912000 $Y=11928000
X6338 24 5807 or03 $T=3019000 11000000 1 180 $X=2968000 $Y=11000000
X6339 24 5808 or03 $T=3019000 11696000 1 180 $X=2968000 $Y=11696000
X6340 24 5809 or03 $T=3019000 11928000 1 180 $X=2968000 $Y=11928000
X6341 24 5810 or03 $T=3075000 11696000 1 180 $X=3024000 $Y=11696000
X6342 24 5811 or03 $T=3075000 11928000 1 180 $X=3024000 $Y=11928000
X6343 24 5812 or03 $T=3131000 11928000 1 180 $X=3080000 $Y=11928000
X6344 24 5813 or03 $T=3187000 11928000 1 180 $X=3136000 $Y=11928000
X6345 24 5814 or03 $T=3512000 12160000 0 0 $X=3512000 $Y=12160000
X6346 24 5815 or03 $T=3712000 13088000 0 0 $X=3712000 $Y=13088000
X6347 24 5816 or03 $T=3808000 13088000 0 0 $X=3808000 $Y=13088000
X6348 24 5817 or03 $T=4048000 12624000 0 0 $X=4048000 $Y=12624000
X6349 24 2316 or03 $T=4048000 13088000 0 0 $X=4048000 $Y=13088000
X6350 24 5818 or03 $T=4088000 13552000 0 0 $X=4088000 $Y=13552000
X6351 24 5819 or03 $T=4104000 12624000 0 0 $X=4104000 $Y=12624000
X6352 24 5820 or03 $T=4136000 13320000 0 0 $X=4136000 $Y=13320000
X6353 24 5821 or03 $T=4184000 13552000 0 0 $X=4184000 $Y=13552000
X6354 24 5822 or03 $T=4443000 12160000 1 180 $X=4392000 $Y=12160000
X6355 24 5823 or03 $T=4499000 12160000 1 180 $X=4448000 $Y=12160000
X6356 24 5824 or03 $T=4888000 13088000 0 0 $X=4888000 $Y=13088000
X6357 24 5825 or03 $T=4960000 12392000 0 0 $X=4960000 $Y=12392000
X6358 24 5826 or03 $T=5035000 13088000 1 180 $X=4984000 $Y=13088000
X6359 24 5827 or03 $T=5091000 13088000 1 180 $X=5040000 $Y=13088000
X6360 24 5828 or03 $T=5120000 12392000 0 0 $X=5120000 $Y=12392000
X6361 24 5829 or03 $T=5120000 12624000 0 0 $X=5120000 $Y=12624000
X6362 24 5830 or03 $T=5227000 12624000 1 180 $X=5176000 $Y=12624000
X6363 24 5831 or03 $T=5339000 12392000 1 180 $X=5288000 $Y=12392000
X6364 24 5832 or03 $T=5379000 12624000 1 180 $X=5328000 $Y=12624000
X6365 24 5833 or03 $T=5395000 13088000 1 180 $X=5344000 $Y=13088000
X6366 24 5834 or03 $T=5483000 13088000 1 180 $X=5432000 $Y=13088000
X6367 24 5835 or03 $T=5539000 13088000 1 180 $X=5488000 $Y=13088000
X6368 24 ICV_36 $T=455000 328000 1 180 $X=392000 $Y=328000
X6369 24 ICV_36 $T=791000 792000 1 180 $X=728000 $Y=792000
X6370 24 ICV_36 $T=919000 1256000 1 180 $X=856000 $Y=1256000
X6371 24 ICV_36 $T=975000 1952000 1 180 $X=912000 $Y=1952000
X6372 24 ICV_36 $T=2327000 1024000 1 180 $X=2264000 $Y=1024000
X6373 24 ICV_36 $T=2687000 2184000 1 180 $X=2624000 $Y=2184000
X6374 24 ICV_36 $T=2695000 1488000 1 180 $X=2632000 $Y=1488000
X6375 24 ICV_36 $T=2895000 1720000 1 180 $X=2832000 $Y=1720000
X6376 24 ICV_36 $T=3551000 96000 1 180 $X=3488000 $Y=96000
X6377 24 ICV_37 $T=375000 2416000 1 180 $X=312000 $Y=2416000
X6378 24 ICV_37 $T=495000 4272000 1 180 $X=432000 $Y=4272000
X6379 24 ICV_37 $T=575000 3344000 1 180 $X=512000 $Y=3344000
X6380 24 ICV_37 $T=951000 2648000 1 180 $X=888000 $Y=2648000
X6381 24 ICV_37 $T=1423000 2880000 1 180 $X=1360000 $Y=2880000
X6382 24 ICV_37 $T=2615000 1952000 1 180 $X=2552000 $Y=1952000
X6383 24 ICV_37 $T=2911000 1488000 1 180 $X=2848000 $Y=1488000
X6384 24 nand03 $T=1185000 2880000 1 180 $X=1144000 $Y=2880000
X6385 24 nand03 $T=1392000 3344000 0 0 $X=1392000 $Y=3344000
X6386 24 nand03 $T=1529000 3344000 1 180 $X=1488000 $Y=3344000
X6387 24 nand03 $T=2248000 1952000 0 0 $X=2248000 $Y=1952000
X6388 24 nand03 $T=2456000 2648000 0 0 $X=2456000 $Y=2648000
X6389 24 nand03 $T=2577000 2648000 1 180 $X=2536000 $Y=2648000
X6390 24 ao32 $T=1616000 3112000 0 0 $X=1616000 $Y=3112000
X6391 24 ao32 $T=2288000 2416000 0 0 $X=2288000 $Y=2416000
X6392 24 ao32 $T=2489500 2416000 1 180 $X=2424000 $Y=2416000
X6393 24 nor02ii $T=441000 8448000 1 180 $X=400000 $Y=8448000
X6394 24 nor02ii $T=481000 8680000 1 180 $X=440000 $Y=8680000
X6395 24 nor02ii $T=528000 8680000 0 0 $X=528000 $Y=8680000
X6396 24 nor02ii $T=617000 8680000 1 180 $X=576000 $Y=8680000
X6397 24 nor02ii $T=841000 8912000 1 180 $X=800000 $Y=8912000
X6398 24 nor02ii $T=889000 8680000 1 180 $X=848000 $Y=8680000
X6399 24 nor02ii $T=889000 8912000 1 180 $X=848000 $Y=8912000
X6400 24 nor02ii $T=1521000 9840000 1 180 $X=1480000 $Y=9840000
X6401 24 nor02ii $T=1569000 9840000 1 180 $X=1528000 $Y=9840000
X6402 24 nor02ii $T=1528000 10072000 0 0 $X=1528000 $Y=10072000
X6403 24 nor02ii $T=1617000 10072000 1 180 $X=1576000 $Y=10072000
X6404 24 nor02ii $T=1632000 1952000 0 0 $X=1632000 $Y=1952000
X6405 24 nor02ii $T=1849000 1952000 1 180 $X=1808000 $Y=1952000
X6406 24 nor02ii $T=2225000 3112000 1 180 $X=2184000 $Y=3112000
X6407 24 nor02ii $T=2408000 3112000 0 0 $X=2408000 $Y=3112000
X6408 24 nand02_2x $T=1921000 2880000 1 180 $X=1888000 $Y=2880000
X6409 24 ICV_38 $T=439000 1256000 1 180 $X=376000 $Y=1256000
X6410 24 ICV_38 $T=511000 3808000 1 180 $X=448000 $Y=3808000
X6411 24 ICV_38 $T=783000 1256000 1 180 $X=720000 $Y=1256000
X6412 24 ICV_38 $T=1887000 792000 1 180 $X=1824000 $Y=792000
X6413 24 ICV_39 $T=375000 2880000 1 180 $X=312000 $Y=2880000
X6414 24 ICV_39 $T=471000 3112000 1 180 $X=408000 $Y=3112000
X6415 24 ICV_39 $T=735000 3576000 1 180 $X=672000 $Y=3576000
X6416 24 ICV_39 $T=1343000 1952000 1 180 $X=1280000 $Y=1952000
X6417 24 ICV_40 $T=504000 560000 0 0 $X=504000 $Y=560000
X6418 24 ICV_40 $T=512000 4040000 0 0 $X=512000 $Y=4040000
X6419 24 ICV_40 $T=624000 3112000 0 0 $X=624000 $Y=3112000
X6420 24 ICV_40 $T=696000 1024000 0 0 $X=696000 $Y=1024000
.ENDS
***************************************
