//
// Verilog description for cell CameraModule, 
// Fri May 12 17:41:22 2017
//
// LeonardoSpectrum Level 3, 2016a.6 
//


module CameraModule ( clk, rst, start, motor_done, nvm_input_address, 
                      nvm_input_data, zero, one, nvm_output_address, 
                      motor_direction, motor_move, done ) ;

    input clk ;
    input rst ;
    input start ;
    input motor_done ;
    input [11:0]nvm_input_address ;
    input [127:0]nvm_input_data ;
    input zero ;
    input one ;
    output [11:0]nvm_output_address ;
    output [0:0]motor_direction ;
    output motor_move ;
    output done ;

    wire ack_from_DMA, write_from_DMA, start_DMA_from_Module, 
         nvm_address_from_Module_11, nvm_address_from_Module_10, 
         nvm_address_from_Module_9, nvm_address_from_Module_8, 
         nvm_address_from_Module_7, nvm_address_from_Module_6, 
         nvm_address_from_Module_5, nvm_address_from_Module_4, 
         nvm_address_from_Module_3, nvm_address_from_Module_2, 
         nvm_address_from_Module_1, nvm_address_from_Module_0, 
         cache_address_from_DMA_7, cache_address_from_DMA_6, 
         cache_address_from_DMA_5, cache_address_from_DMA_4, 
         cache_address_from_DMA_3, cache_address_from_DMA_2, 
         cache_address_from_DMA_1, cache_address_from_DMA_0, 
         cache_address_from_Module_7, cache_address_from_Module_6, 
         cache_address_from_Module_5, cache_address_from_Module_4, 
         cache_address_from_Module_3, cache_address_from_Module_2, 
         cache_address_from_Module_1, cache_address_from_Module_0, 
         address_to_cache_7, address_to_cache_6, address_to_cache_5, 
         address_to_cache_4, address_to_cache_3, address_to_cache_2, 
         address_to_cache_1, address_to_cache_0, data_from_DMA_7, 
         data_from_DMA_6, data_from_DMA_5, data_from_DMA_4, data_from_DMA_3, 
         data_from_DMA_2, data_from_DMA_1, data_from_DMA_0, data_from_cache_7, 
         data_from_cache_6, data_from_cache_5, data_from_cache_4, 
         data_from_cache_3, data_from_cache_2, data_from_cache_1, 
         data_from_cache_0, nx241, nx247, nx249;
    wire [4:0] \$dummy ;




    nbit_mux2x1_8 mux (.input1 ({cache_address_from_Module_7,
                  cache_address_from_Module_6,cache_address_from_Module_5,
                  cache_address_from_Module_4,cache_address_from_Module_3,
                  cache_address_from_Module_2,cache_address_from_Module_1,
                  cache_address_from_Module_0}), .input2 ({
                  cache_address_from_DMA_7,cache_address_from_DMA_6,
                  cache_address_from_DMA_5,cache_address_from_DMA_4,
                  cache_address_from_DMA_3,cache_address_from_DMA_2,
                  cache_address_from_DMA_1,cache_address_from_DMA_0}), .s0 (
                  nx247), .\output  ({address_to_cache_7,address_to_cache_6,
                  address_to_cache_5,address_to_cache_4,address_to_cache_3,
                  address_to_cache_2,address_to_cache_1,address_to_cache_0})) ;
    CacheMemory cache (.clk (clk), .rst (rst), .write_en (nx249), .address ({
                address_to_cache_7,address_to_cache_6,address_to_cache_5,
                address_to_cache_4,address_to_cache_3,address_to_cache_2,
                address_to_cache_1,address_to_cache_0}), .datain ({
                data_from_DMA_7,data_from_DMA_6,data_from_DMA_5,data_from_DMA_4,
                data_from_DMA_3,data_from_DMA_2,data_from_DMA_1,data_from_DMA_0}
                ), .dataout ({data_from_cache_7,data_from_cache_6,
                data_from_cache_5,data_from_cache_4,data_from_cache_3,
                data_from_cache_2,data_from_cache_1,data_from_cache_0})) ;
    \module  algo_module (.clk (clk), .rst (rst), .ack (ack_from_DMA), .start (
             start), .move_done (motor_done), .nvm_address_in ({
             nvm_input_address[11],nvm_input_address[10],nvm_input_address[9],
             nvm_input_address[8],nvm_input_address[7],nvm_input_address[6],
             nvm_input_address[5],nvm_input_address[4],nvm_input_address[3],
             nvm_input_address[2],nvm_input_address[1],nvm_input_address[0]}), .cache_data_in (
             {data_from_cache_7,data_from_cache_6,data_from_cache_5,
             data_from_cache_4,data_from_cache_3,data_from_cache_2,
             data_from_cache_1,data_from_cache_0}), .zero (zero), .one (one), .cache_address_out (
             {cache_address_from_Module_7,cache_address_from_Module_6,
             cache_address_from_Module_5,cache_address_from_Module_4,
             cache_address_from_Module_3,cache_address_from_Module_2,
             cache_address_from_Module_1,cache_address_from_Module_0}), .move (
             motor_move), .start_dma (start_DMA_from_Module), .done (done), .direction (
             {motor_direction[0]}), .nvm_address_out ({
             nvm_address_from_Module_11,nvm_address_from_Module_10,
             nvm_address_from_Module_9,nvm_address_from_Module_8,
             nvm_address_from_Module_7,nvm_address_from_Module_6,
             nvm_address_from_Module_5,nvm_address_from_Module_4,
             nvm_address_from_Module_3,nvm_address_from_Module_2,
             nvm_address_from_Module_1,nvm_address_from_Module_0}), .state_out (
             {\$dummy [0],\$dummy [1],\$dummy [2],\$dummy [3],\$dummy [4]})) ;
    DMA DMA_module (.clk (clk), .rst (rst), .start_DMA (nx241), .Data_in ({
        nvm_input_data[127],nvm_input_data[126],nvm_input_data[125],
        nvm_input_data[124],nvm_input_data[123],nvm_input_data[122],
        nvm_input_data[121],nvm_input_data[120],nvm_input_data[119],
        nvm_input_data[118],nvm_input_data[117],nvm_input_data[116],
        nvm_input_data[115],nvm_input_data[114],nvm_input_data[113],
        nvm_input_data[112],nvm_input_data[111],nvm_input_data[110],
        nvm_input_data[109],nvm_input_data[108],nvm_input_data[107],
        nvm_input_data[106],nvm_input_data[105],nvm_input_data[104],
        nvm_input_data[103],nvm_input_data[102],nvm_input_data[101],
        nvm_input_data[100],nvm_input_data[99],nvm_input_data[98],
        nvm_input_data[97],nvm_input_data[96],nvm_input_data[95],
        nvm_input_data[94],nvm_input_data[93],nvm_input_data[92],
        nvm_input_data[91],nvm_input_data[90],nvm_input_data[89],
        nvm_input_data[88],nvm_input_data[87],nvm_input_data[86],
        nvm_input_data[85],nvm_input_data[84],nvm_input_data[83],
        nvm_input_data[82],nvm_input_data[81],nvm_input_data[80],
        nvm_input_data[79],nvm_input_data[78],nvm_input_data[77],
        nvm_input_data[76],nvm_input_data[75],nvm_input_data[74],
        nvm_input_data[73],nvm_input_data[72],nvm_input_data[71],
        nvm_input_data[70],nvm_input_data[69],nvm_input_data[68],
        nvm_input_data[67],nvm_input_data[66],nvm_input_data[65],
        nvm_input_data[64],nvm_input_data[63],nvm_input_data[62],
        nvm_input_data[61],nvm_input_data[60],nvm_input_data[59],
        nvm_input_data[58],nvm_input_data[57],nvm_input_data[56],
        nvm_input_data[55],nvm_input_data[54],nvm_input_data[53],
        nvm_input_data[52],nvm_input_data[51],nvm_input_data[50],
        nvm_input_data[49],nvm_input_data[48],nvm_input_data[47],
        nvm_input_data[46],nvm_input_data[45],nvm_input_data[44],
        nvm_input_data[43],nvm_input_data[42],nvm_input_data[41],
        nvm_input_data[40],nvm_input_data[39],nvm_input_data[38],
        nvm_input_data[37],nvm_input_data[36],nvm_input_data[35],
        nvm_input_data[34],nvm_input_data[33],nvm_input_data[32],
        nvm_input_data[31],nvm_input_data[30],nvm_input_data[29],
        nvm_input_data[28],nvm_input_data[27],nvm_input_data[26],
        nvm_input_data[25],nvm_input_data[24],nvm_input_data[23],
        nvm_input_data[22],nvm_input_data[21],nvm_input_data[20],
        nvm_input_data[19],nvm_input_data[18],nvm_input_data[17],
        nvm_input_data[16],nvm_input_data[15],nvm_input_data[14],
        nvm_input_data[13],nvm_input_data[12],nvm_input_data[11],
        nvm_input_data[10],nvm_input_data[9],nvm_input_data[8],nvm_input_data[7]
        ,nvm_input_data[6],nvm_input_data[5],nvm_input_data[4],nvm_input_data[3]
        ,nvm_input_data[2],nvm_input_data[1],nvm_input_data[0]}), .NVM_addr_in (
        {nvm_address_from_Module_11,nvm_address_from_Module_10,
        nvm_address_from_Module_9,nvm_address_from_Module_8,
        nvm_address_from_Module_7,nvm_address_from_Module_6,
        nvm_address_from_Module_5,nvm_address_from_Module_4,
        nvm_address_from_Module_3,nvm_address_from_Module_2,
        nvm_address_from_Module_1,nvm_address_from_Module_0}), .zero (zero), .one (
        one), .write_signal (write_from_DMA), .Ack (ack_from_DMA), .Data_out ({
        data_from_DMA_7,data_from_DMA_6,data_from_DMA_5,data_from_DMA_4,
        data_from_DMA_3,data_from_DMA_2,data_from_DMA_1,data_from_DMA_0}), .cache_addr (
        {cache_address_from_DMA_7,cache_address_from_DMA_6,
        cache_address_from_DMA_5,cache_address_from_DMA_4,
        cache_address_from_DMA_3,cache_address_from_DMA_2,
        cache_address_from_DMA_1,cache_address_from_DMA_0}), .NVM_addr_out ({
        nvm_output_address[11],nvm_output_address[10],nvm_output_address[9],
        nvm_output_address[8],nvm_output_address[7],nvm_output_address[6],
        nvm_output_address[5],nvm_output_address[4],nvm_output_address[3],
        nvm_output_address[2],nvm_output_address[1],nvm_output_address[0]})) ;
    buf02 ix240 (.Y (nx241), .A (start_DMA_from_Module)) ;
    buf02 ix246 (.Y (nx247), .A (write_from_DMA)) ;
    buf02 ix248 (.Y (nx249), .A (write_from_DMA)) ;
endmodule


module DMA ( clk, rst, start_DMA, Data_in, NVM_addr_in, zero, one, write_signal, 
             Ack, Data_out, cache_addr, NVM_addr_out ) ;

    input clk ;
    input rst ;
    input start_DMA ;
    input [127:0]Data_in ;
    input [11:0]NVM_addr_in ;
    input zero ;
    input one ;
    output write_signal ;
    output Ack ;
    output [7:0]Data_out ;
    output [7:0]cache_addr ;
    output [11:0]NVM_addr_out ;

    wire cache_adder_out_7, cache_adder_out_6, cache_adder_out_5, 
         cache_adder_out_4, cache_adder_out_3, cache_adder_out_2, 
         cache_adder_out_1, cache_adder_out_0, NVM_adder_out_11, 
         NVM_adder_out_10, NVM_adder_out_9, NVM_adder_out_8, NVM_adder_out_7, 
         NVM_adder_out_6, NVM_adder_out_5, NVM_adder_out_4, NVM_adder_out_3, 
         NVM_adder_out_2, NVM_adder_out_1, NVM_adder_out_0, 
         NVM_address_Mux_out_11, NVM_address_Mux_out_10, NVM_address_Mux_out_9, 
         NVM_address_Mux_out_8, NVM_address_Mux_out_7, NVM_address_Mux_out_6, 
         NVM_address_Mux_out_5, NVM_address_Mux_out_4, NVM_address_Mux_out_3, 
         NVM_address_Mux_out_2, NVM_address_Mux_out_1, NVM_address_Mux_out_0, 
         row_done, rows_done, signals_4, signals_3, signals_1;
    wire [0:0] \$dummy ;




    DMACU controlUnit (.clk (clk), .reset (rst), .start_DMA (start_DMA), .Rows_Done (
          rows_done), .Row_Done (row_done), .signals ({write_signal,signals_4,
          signals_3,\$dummy [0],signals_1,Ack})) ;
    nbit_Register_8 R_Cache_addr (.Clk (clk), .rst (signals_1), .enable (
                    write_signal), .d ({cache_adder_out_7,cache_adder_out_6,
                    cache_adder_out_5,cache_adder_out_4,cache_adder_out_3,
                    cache_adder_out_2,cache_adder_out_1,cache_adder_out_0}), .rst_value (
                    {zero,zero,zero,zero,zero,zero,zero,zero}), .q ({
                    cache_addr[7],cache_addr[6],cache_addr[5],cache_addr[4],
                    cache_addr[3],cache_addr[2],cache_addr[1],cache_addr[0]})) ;
    nbit_Register_12 R_NVM_addr (.Clk (clk), .rst (signals_1), .enable (
                     signals_3), .d ({NVM_address_Mux_out_11,
                     NVM_address_Mux_out_10,NVM_address_Mux_out_9,
                     NVM_address_Mux_out_8,NVM_address_Mux_out_7,
                     NVM_address_Mux_out_6,NVM_address_Mux_out_5,
                     NVM_address_Mux_out_4,NVM_address_Mux_out_3,
                     NVM_address_Mux_out_2,NVM_address_Mux_out_1,
                     NVM_address_Mux_out_0}), .rst_value ({zero,zero,zero,zero,
                     zero,zero,zero,zero,zero,zero,zero,zero}), .q ({
                     NVM_addr_out[11],NVM_addr_out[10],NVM_addr_out[9],
                     NVM_addr_out[8],NVM_addr_out[7],NVM_addr_out[6],
                     NVM_addr_out[5],NVM_addr_out[4],NVM_addr_out[3],
                     NVM_addr_out[2],NVM_addr_out[1],NVM_addr_out[0]})) ;
    nbit_adder_8 u1 (.a ({cache_addr[7],cache_addr[6],cache_addr[5],
                 cache_addr[4],cache_addr[3],cache_addr[2],cache_addr[1],
                 cache_addr[0]}), .b ({zero,zero,zero,zero,zero,zero,zero,zero})
                 , .cin (one), .add_out ({cache_adder_out_7,cache_adder_out_6,
                 cache_adder_out_5,cache_adder_out_4,cache_adder_out_3,
                 cache_adder_out_2,cache_adder_out_1,cache_adder_out_0})) ;
    nbit_adder_12 u2 (.a ({NVM_addr_out[11],NVM_addr_out[10],NVM_addr_out[9],
                  NVM_addr_out[8],NVM_addr_out[7],NVM_addr_out[6],
                  NVM_addr_out[5],NVM_addr_out[4],NVM_addr_out[3],
                  NVM_addr_out[2],NVM_addr_out[1],NVM_addr_out[0]}), .b ({zero,
                  zero,zero,zero,zero,zero,zero,one,zero,zero,zero,zero}), .cin (
                  zero), .add_out ({NVM_adder_out_11,NVM_adder_out_10,
                  NVM_adder_out_9,NVM_adder_out_8,NVM_adder_out_7,
                  NVM_adder_out_6,NVM_adder_out_5,NVM_adder_out_4,
                  NVM_adder_out_3,NVM_adder_out_2,NVM_adder_out_1,
                  NVM_adder_out_0})) ;
    mux16x1 u3 (.x0 ({Data_in[127],Data_in[126],Data_in[125],Data_in[124],
            Data_in[123],Data_in[122],Data_in[121],Data_in[120]}), .x1 ({
            Data_in[119],Data_in[118],Data_in[117],Data_in[116],Data_in[115],
            Data_in[114],Data_in[113],Data_in[112]}), .x2 ({Data_in[111],
            Data_in[110],Data_in[109],Data_in[108],Data_in[107],Data_in[106],
            Data_in[105],Data_in[104]}), .x3 ({Data_in[103],Data_in[102],
            Data_in[101],Data_in[100],Data_in[99],Data_in[98],Data_in[97],
            Data_in[96]}), .x4 ({Data_in[95],Data_in[94],Data_in[93],Data_in[92]
            ,Data_in[91],Data_in[90],Data_in[89],Data_in[88]}), .x5 ({
            Data_in[87],Data_in[86],Data_in[85],Data_in[84],Data_in[83],
            Data_in[82],Data_in[81],Data_in[80]}), .x6 ({Data_in[79],Data_in[78]
            ,Data_in[77],Data_in[76],Data_in[75],Data_in[74],Data_in[73],
            Data_in[72]}), .x7 ({Data_in[71],Data_in[70],Data_in[69],Data_in[68]
            ,Data_in[67],Data_in[66],Data_in[65],Data_in[64]}), .x8 ({
            Data_in[63],Data_in[62],Data_in[61],Data_in[60],Data_in[59],
            Data_in[58],Data_in[57],Data_in[56]}), .x9 ({Data_in[55],Data_in[54]
            ,Data_in[53],Data_in[52],Data_in[51],Data_in[50],Data_in[49],
            Data_in[48]}), .x10 ({Data_in[47],Data_in[46],Data_in[45],
            Data_in[44],Data_in[43],Data_in[42],Data_in[41],Data_in[40]}), .x11 (
            {Data_in[39],Data_in[38],Data_in[37],Data_in[36],Data_in[35],
            Data_in[34],Data_in[33],Data_in[32]}), .x12 ({Data_in[31],
            Data_in[30],Data_in[29],Data_in[28],Data_in[27],Data_in[26],
            Data_in[25],Data_in[24]}), .x13 ({Data_in[23],Data_in[22],
            Data_in[21],Data_in[20],Data_in[19],Data_in[18],Data_in[17],
            Data_in[16]}), .x14 ({Data_in[15],Data_in[14],Data_in[13],
            Data_in[12],Data_in[11],Data_in[10],Data_in[9],Data_in[8]}), .x15 ({
            Data_in[7],Data_in[6],Data_in[5],Data_in[4],Data_in[3],Data_in[2],
            Data_in[1],Data_in[0]}), .sel ({cache_addr[3],cache_addr[2],
            cache_addr[1],cache_addr[0]}), .y ({Data_out[7],Data_out[6],
            Data_out[5],Data_out[4],Data_out[3],Data_out[2],Data_out[1],
            Data_out[0]})) ;
    nbit_mux2x1_12 u4 (.input1 ({NVM_adder_out_11,NVM_adder_out_10,
                   NVM_adder_out_9,NVM_adder_out_8,NVM_adder_out_7,
                   NVM_adder_out_6,NVM_adder_out_5,NVM_adder_out_4,
                   NVM_adder_out_3,NVM_adder_out_2,NVM_adder_out_1,
                   NVM_adder_out_0}), .input2 ({NVM_addr_in[11],NVM_addr_in[10],
                   NVM_addr_in[9],NVM_addr_in[8],NVM_addr_in[7],NVM_addr_in[6],
                   NVM_addr_in[5],NVM_addr_in[4],NVM_addr_in[3],NVM_addr_in[2],
                   NVM_addr_in[1],NVM_addr_in[0]}), .s0 (signals_4), .\output  (
                   {NVM_address_Mux_out_11,NVM_address_Mux_out_10,
                   NVM_address_Mux_out_9,NVM_address_Mux_out_8,
                   NVM_address_Mux_out_7,NVM_address_Mux_out_6,
                   NVM_address_Mux_out_5,NVM_address_Mux_out_4,
                   NVM_address_Mux_out_3,NVM_address_Mux_out_2,
                   NVM_address_Mux_out_1,NVM_address_Mux_out_0})) ;
    and04 ix5 (.Y (rows_done), .A0 (cache_addr[7]), .A1 (cache_addr[6]), .A2 (
          cache_addr[5]), .A3 (cache_addr[4])) ;
    and04 ix11 (.Y (row_done), .A0 (cache_addr[3]), .A1 (cache_addr[2]), .A2 (
          cache_addr[1]), .A3 (cache_addr[0])) ;
endmodule


module nbit_mux2x1_12 ( input1, input2, s0, \output  ) ;

    input [11:0]input1 ;
    input [11:0]input2 ;
    input s0 ;
    output [11:0]\output  ;

    wire nx185, nx187;



    mux21_ni ix7 (.Y (\output [0]), .A0 (input1[0]), .A1 (input2[0]), .S0 (nx185
             )) ;
    mux21_ni ix15 (.Y (\output [1]), .A0 (input1[1]), .A1 (input2[1]), .S0 (
             nx185)) ;
    mux21_ni ix23 (.Y (\output [2]), .A0 (input1[2]), .A1 (input2[2]), .S0 (
             nx185)) ;
    mux21_ni ix31 (.Y (\output [3]), .A0 (input1[3]), .A1 (input2[3]), .S0 (
             nx185)) ;
    mux21_ni ix39 (.Y (\output [4]), .A0 (input1[4]), .A1 (input2[4]), .S0 (
             nx185)) ;
    mux21_ni ix47 (.Y (\output [5]), .A0 (input1[5]), .A1 (input2[5]), .S0 (
             nx185)) ;
    mux21_ni ix55 (.Y (\output [6]), .A0 (input1[6]), .A1 (input2[6]), .S0 (
             nx185)) ;
    mux21_ni ix63 (.Y (\output [7]), .A0 (input1[7]), .A1 (input2[7]), .S0 (
             nx187)) ;
    mux21_ni ix71 (.Y (\output [8]), .A0 (input1[8]), .A1 (input2[8]), .S0 (
             nx187)) ;
    mux21_ni ix79 (.Y (\output [9]), .A0 (input1[9]), .A1 (input2[9]), .S0 (
             nx187)) ;
    mux21_ni ix87 (.Y (\output [10]), .A0 (input1[10]), .A1 (input2[10]), .S0 (
             nx187)) ;
    mux21_ni ix95 (.Y (\output [11]), .A0 (input1[11]), .A1 (input2[11]), .S0 (
             nx187)) ;
    buf02 ix184 (.Y (nx185), .A (s0)) ;
    buf02 ix186 (.Y (nx187), .A (s0)) ;
endmodule


module mux16x1 ( x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, 
                 x15, sel, y ) ;

    input [7:0]x0 ;
    input [7:0]x1 ;
    input [7:0]x2 ;
    input [7:0]x3 ;
    input [7:0]x4 ;
    input [7:0]x5 ;
    input [7:0]x6 ;
    input [7:0]x7 ;
    input [7:0]x8 ;
    input [7:0]x9 ;
    input [7:0]x10 ;
    input [7:0]x11 ;
    input [7:0]x12 ;
    input [7:0]x13 ;
    input [7:0]x14 ;
    input [7:0]x15 ;
    input [3:0]sel ;
    output [7:0]y ;

    wire nx10, nx18, nx32, nx36, nx48, nx54, nx60, nx68, nx76, nx78, nx82, nx88, 
         nx92, nx100, nx104, nx110, nx114, nx122, nx154, nx184, nx216, nx246, 
         nx278, nx308, nx340, nx370, nx402, nx432, nx464, nx494, nx526, nx556, 
         nx255, nx259, nx261, nx265, nx267, nx271, nx273, nx277, nx279, nx281, 
         nx285, nx289, nx293, nx295, nx301, nx307, nx313, nx319, nx329, nx331, 
         nx333, nx335, nx339, nx341, nx343, nx345, nx351, nx353, nx355, nx357, 
         nx361, nx363, nx365, nx367, nx373, nx375, nx377, nx379, nx383, nx385, 
         nx387, nx389, nx395, nx397, nx399, nx401, nx405, nx407, nx409, nx411, 
         nx417, nx419, nx421, nx423, nx427, nx429, nx431, nx433, nx439, nx441, 
         nx443, nx445, nx449, nx451, nx453, nx455, nx461, nx463, nx465, nx467, 
         nx471, nx473, nx475, nx477, nx484, nx486, nx492, nx495, nx497, nx499;



    or02 ix125 (.Y (y[0]), .A0 (nx122), .A1 (nx76)) ;
    nand04 ix123 (.Y (nx122), .A0 (nx255), .A1 (nx267), .A2 (nx281), .A3 (nx289)
           ) ;
    aoi22 ix256 (.Y (nx255), .A0 (x4[0]), .A1 (nx114), .B0 (x7[0]), .B1 (nx110)
          ) ;
    nor03_2x ix115 (.Y (nx114), .A0 (nx497), .A1 (nx499), .A2 (nx259)) ;
    nand02 ix260 (.Y (nx259), .A0 (nx261), .A1 (nx495)) ;
    inv01 ix262 (.Y (nx261), .A (sel[3])) ;
    nor02_2x ix111 (.Y (nx110), .A0 (nx265), .A1 (nx259)) ;
    nand02 ix266 (.Y (nx265), .A0 (nx497), .A1 (nx499)) ;
    aoi22 ix268 (.Y (nx267), .A0 (x11[0]), .A1 (nx100), .B0 (x6[0]), .B1 (nx104)
          ) ;
    nor02_2x ix104 (.Y (nx100), .A0 (nx265), .A1 (nx271)) ;
    nand02 ix272 (.Y (nx271), .A0 (nx492), .A1 (nx273)) ;
    inv01 ix274 (.Y (nx273), .A (sel[2])) ;
    nor02_2x ix106 (.Y (nx104), .A0 (nx277), .A1 (nx259)) ;
    nand02 ix278 (.Y (nx277), .A0 (nx497), .A1 (nx279)) ;
    inv01 ix280 (.Y (nx279), .A (sel[0])) ;
    aoi22 ix282 (.Y (nx281), .A0 (x15[0]), .A1 (nx88), .B0 (x12[0]), .B1 (nx92)
          ) ;
    nor02_2x ix89 (.Y (nx88), .A0 (nx285), .A1 (nx265)) ;
    nand02 ix286 (.Y (nx285), .A0 (nx492), .A1 (nx495)) ;
    nor03_2x ix93 (.Y (nx92), .A0 (nx285), .A1 (nx497), .A2 (nx499)) ;
    aoi22 ix290 (.Y (nx289), .A0 (x1[0]), .A1 (nx82), .B0 (x0[0]), .B1 (nx484)
          ) ;
    nor03_2x ix83 (.Y (nx82), .A0 (nx492), .A1 (nx495), .A2 (nx293)) ;
    nand02 ix294 (.Y (nx293), .A0 (nx295), .A1 (nx499)) ;
    inv01 ix296 (.Y (nx295), .A (sel[1])) ;
    nor04 ix79 (.Y (nx78), .A0 (nx497), .A1 (nx499), .A2 (nx492), .A3 (nx495)) ;
    nand04 ix77 (.Y (nx76), .A0 (nx301), .A1 (nx307), .A2 (nx313), .A3 (nx319)
           ) ;
    aoi22 ix302 (.Y (nx301), .A0 (x5[0]), .A1 (nx68), .B0 (x14[0]), .B1 (nx60)
          ) ;
    nor02_2x ix69 (.Y (nx68), .A0 (nx259), .A1 (nx293)) ;
    nor02_2x ix61 (.Y (nx60), .A0 (nx285), .A1 (nx277)) ;
    aoi22 ix308 (.Y (nx307), .A0 (x13[0]), .A1 (nx54), .B0 (x9[0]), .B1 (nx48)
          ) ;
    nor02_2x ix55 (.Y (nx54), .A0 (nx285), .A1 (nx293)) ;
    nor02_2x ix49 (.Y (nx48), .A0 (nx271), .A1 (nx293)) ;
    aoi22 ix314 (.Y (nx313), .A0 (x3[0]), .A1 (nx32), .B0 (x2[0]), .B1 (nx36)) ;
    nor03_2x ix33 (.Y (nx32), .A0 (nx265), .A1 (nx492), .A2 (nx495)) ;
    nor03_2x ix37 (.Y (nx36), .A0 (nx277), .A1 (nx492), .A2 (nx495)) ;
    aoi22 ix320 (.Y (nx319), .A0 (x8[0]), .A1 (nx10), .B0 (x10[0]), .B1 (nx18)
          ) ;
    nor03_2x ix11 (.Y (nx10), .A0 (nx497), .A1 (nx499), .A2 (nx271)) ;
    nor02_2x ix19 (.Y (nx18), .A0 (nx277), .A1 (nx271)) ;
    or02 ix187 (.Y (y[1]), .A0 (nx184), .A1 (nx154)) ;
    nand04 ix185 (.Y (nx184), .A0 (nx329), .A1 (nx331), .A2 (nx333), .A3 (nx335)
           ) ;
    aoi22 ix330 (.Y (nx329), .A0 (x4[1]), .A1 (nx114), .B0 (x7[1]), .B1 (nx110)
          ) ;
    aoi22 ix332 (.Y (nx331), .A0 (x11[1]), .A1 (nx100), .B0 (x6[1]), .B1 (nx104)
          ) ;
    aoi22 ix334 (.Y (nx333), .A0 (x15[1]), .A1 (nx88), .B0 (x12[1]), .B1 (nx92)
          ) ;
    aoi22 ix336 (.Y (nx335), .A0 (x1[1]), .A1 (nx82), .B0 (x0[1]), .B1 (nx484)
          ) ;
    nand04 ix155 (.Y (nx154), .A0 (nx339), .A1 (nx341), .A2 (nx343), .A3 (nx345)
           ) ;
    aoi22 ix340 (.Y (nx339), .A0 (x5[1]), .A1 (nx68), .B0 (x14[1]), .B1 (nx60)
          ) ;
    aoi22 ix342 (.Y (nx341), .A0 (x13[1]), .A1 (nx54), .B0 (x9[1]), .B1 (nx48)
          ) ;
    aoi22 ix344 (.Y (nx343), .A0 (x3[1]), .A1 (nx32), .B0 (x2[1]), .B1 (nx36)) ;
    aoi22 ix346 (.Y (nx345), .A0 (x8[1]), .A1 (nx10), .B0 (x10[1]), .B1 (nx18)
          ) ;
    or02 ix249 (.Y (y[2]), .A0 (nx246), .A1 (nx216)) ;
    nand04 ix247 (.Y (nx246), .A0 (nx351), .A1 (nx353), .A2 (nx355), .A3 (nx357)
           ) ;
    aoi22 ix352 (.Y (nx351), .A0 (x4[2]), .A1 (nx114), .B0 (x7[2]), .B1 (nx110)
          ) ;
    aoi22 ix354 (.Y (nx353), .A0 (x11[2]), .A1 (nx100), .B0 (x6[2]), .B1 (nx104)
          ) ;
    aoi22 ix356 (.Y (nx355), .A0 (x15[2]), .A1 (nx88), .B0 (x12[2]), .B1 (nx92)
          ) ;
    aoi22 ix358 (.Y (nx357), .A0 (x1[2]), .A1 (nx82), .B0 (x0[2]), .B1 (nx484)
          ) ;
    nand04 ix217 (.Y (nx216), .A0 (nx361), .A1 (nx363), .A2 (nx365), .A3 (nx367)
           ) ;
    aoi22 ix362 (.Y (nx361), .A0 (x5[2]), .A1 (nx68), .B0 (x14[2]), .B1 (nx60)
          ) ;
    aoi22 ix364 (.Y (nx363), .A0 (x13[2]), .A1 (nx54), .B0 (x9[2]), .B1 (nx48)
          ) ;
    aoi22 ix366 (.Y (nx365), .A0 (x3[2]), .A1 (nx32), .B0 (x2[2]), .B1 (nx36)) ;
    aoi22 ix368 (.Y (nx367), .A0 (x8[2]), .A1 (nx10), .B0 (x10[2]), .B1 (nx18)
          ) ;
    or02 ix311 (.Y (y[3]), .A0 (nx308), .A1 (nx278)) ;
    nand04 ix309 (.Y (nx308), .A0 (nx373), .A1 (nx375), .A2 (nx377), .A3 (nx379)
           ) ;
    aoi22 ix374 (.Y (nx373), .A0 (x4[3]), .A1 (nx114), .B0 (x7[3]), .B1 (nx110)
          ) ;
    aoi22 ix376 (.Y (nx375), .A0 (x11[3]), .A1 (nx100), .B0 (x6[3]), .B1 (nx104)
          ) ;
    aoi22 ix378 (.Y (nx377), .A0 (x15[3]), .A1 (nx88), .B0 (x12[3]), .B1 (nx92)
          ) ;
    aoi22 ix380 (.Y (nx379), .A0 (x1[3]), .A1 (nx82), .B0 (x0[3]), .B1 (nx484)
          ) ;
    nand04 ix279 (.Y (nx278), .A0 (nx383), .A1 (nx385), .A2 (nx387), .A3 (nx389)
           ) ;
    aoi22 ix384 (.Y (nx383), .A0 (x5[3]), .A1 (nx68), .B0 (x14[3]), .B1 (nx60)
          ) ;
    aoi22 ix386 (.Y (nx385), .A0 (x13[3]), .A1 (nx54), .B0 (x9[3]), .B1 (nx48)
          ) ;
    aoi22 ix388 (.Y (nx387), .A0 (x3[3]), .A1 (nx32), .B0 (x2[3]), .B1 (nx36)) ;
    aoi22 ix390 (.Y (nx389), .A0 (x8[3]), .A1 (nx10), .B0 (x10[3]), .B1 (nx18)
          ) ;
    or02 ix373 (.Y (y[4]), .A0 (nx370), .A1 (nx340)) ;
    nand04 ix371 (.Y (nx370), .A0 (nx395), .A1 (nx397), .A2 (nx399), .A3 (nx401)
           ) ;
    aoi22 ix396 (.Y (nx395), .A0 (x4[4]), .A1 (nx114), .B0 (x7[4]), .B1 (nx110)
          ) ;
    aoi22 ix398 (.Y (nx397), .A0 (x11[4]), .A1 (nx100), .B0 (x6[4]), .B1 (nx104)
          ) ;
    aoi22 ix400 (.Y (nx399), .A0 (x15[4]), .A1 (nx88), .B0 (x12[4]), .B1 (nx92)
          ) ;
    aoi22 ix402 (.Y (nx401), .A0 (x1[4]), .A1 (nx82), .B0 (x0[4]), .B1 (nx484)
          ) ;
    nand04 ix341 (.Y (nx340), .A0 (nx405), .A1 (nx407), .A2 (nx409), .A3 (nx411)
           ) ;
    aoi22 ix406 (.Y (nx405), .A0 (x5[4]), .A1 (nx68), .B0 (x14[4]), .B1 (nx60)
          ) ;
    aoi22 ix408 (.Y (nx407), .A0 (x13[4]), .A1 (nx54), .B0 (x9[4]), .B1 (nx48)
          ) ;
    aoi22 ix410 (.Y (nx409), .A0 (x3[4]), .A1 (nx32), .B0 (x2[4]), .B1 (nx36)) ;
    aoi22 ix412 (.Y (nx411), .A0 (x8[4]), .A1 (nx10), .B0 (x10[4]), .B1 (nx18)
          ) ;
    or02 ix435 (.Y (y[5]), .A0 (nx432), .A1 (nx402)) ;
    nand04 ix433 (.Y (nx432), .A0 (nx417), .A1 (nx419), .A2 (nx421), .A3 (nx423)
           ) ;
    aoi22 ix418 (.Y (nx417), .A0 (x4[5]), .A1 (nx114), .B0 (x7[5]), .B1 (nx110)
          ) ;
    aoi22 ix420 (.Y (nx419), .A0 (x11[5]), .A1 (nx100), .B0 (x6[5]), .B1 (nx104)
          ) ;
    aoi22 ix422 (.Y (nx421), .A0 (x15[5]), .A1 (nx88), .B0 (x12[5]), .B1 (nx92)
          ) ;
    aoi22 ix424 (.Y (nx423), .A0 (x1[5]), .A1 (nx82), .B0 (x0[5]), .B1 (nx484)
          ) ;
    nand04 ix403 (.Y (nx402), .A0 (nx427), .A1 (nx429), .A2 (nx431), .A3 (nx433)
           ) ;
    aoi22 ix428 (.Y (nx427), .A0 (x5[5]), .A1 (nx68), .B0 (x14[5]), .B1 (nx60)
          ) ;
    aoi22 ix430 (.Y (nx429), .A0 (x13[5]), .A1 (nx54), .B0 (x9[5]), .B1 (nx48)
          ) ;
    aoi22 ix432 (.Y (nx431), .A0 (x3[5]), .A1 (nx32), .B0 (x2[5]), .B1 (nx36)) ;
    aoi22 ix434 (.Y (nx433), .A0 (x8[5]), .A1 (nx10), .B0 (x10[5]), .B1 (nx18)
          ) ;
    or02 ix497 (.Y (y[6]), .A0 (nx494), .A1 (nx464)) ;
    nand04 ix495 (.Y (nx494), .A0 (nx439), .A1 (nx441), .A2 (nx443), .A3 (nx445)
           ) ;
    aoi22 ix440 (.Y (nx439), .A0 (x4[6]), .A1 (nx114), .B0 (x7[6]), .B1 (nx110)
          ) ;
    aoi22 ix442 (.Y (nx441), .A0 (x11[6]), .A1 (nx100), .B0 (x6[6]), .B1 (nx104)
          ) ;
    aoi22 ix444 (.Y (nx443), .A0 (x15[6]), .A1 (nx88), .B0 (x12[6]), .B1 (nx92)
          ) ;
    aoi22 ix446 (.Y (nx445), .A0 (x1[6]), .A1 (nx82), .B0 (x0[6]), .B1 (nx484)
          ) ;
    nand04 ix465 (.Y (nx464), .A0 (nx449), .A1 (nx451), .A2 (nx453), .A3 (nx455)
           ) ;
    aoi22 ix450 (.Y (nx449), .A0 (x5[6]), .A1 (nx68), .B0 (x14[6]), .B1 (nx60)
          ) ;
    aoi22 ix452 (.Y (nx451), .A0 (x13[6]), .A1 (nx54), .B0 (x9[6]), .B1 (nx48)
          ) ;
    aoi22 ix454 (.Y (nx453), .A0 (x3[6]), .A1 (nx32), .B0 (x2[6]), .B1 (nx36)) ;
    aoi22 ix456 (.Y (nx455), .A0 (x8[6]), .A1 (nx10), .B0 (x10[6]), .B1 (nx18)
          ) ;
    or02 ix559 (.Y (y[7]), .A0 (nx556), .A1 (nx526)) ;
    nand04 ix557 (.Y (nx556), .A0 (nx461), .A1 (nx463), .A2 (nx465), .A3 (nx467)
           ) ;
    aoi22 ix462 (.Y (nx461), .A0 (x4[7]), .A1 (nx114), .B0 (x7[7]), .B1 (nx110)
          ) ;
    aoi22 ix464 (.Y (nx463), .A0 (x11[7]), .A1 (nx100), .B0 (x6[7]), .B1 (nx104)
          ) ;
    aoi22 ix466 (.Y (nx465), .A0 (x15[7]), .A1 (nx88), .B0 (x12[7]), .B1 (nx92)
          ) ;
    aoi22 ix468 (.Y (nx467), .A0 (x1[7]), .A1 (nx82), .B0 (x0[7]), .B1 (nx486)
          ) ;
    nand04 ix527 (.Y (nx526), .A0 (nx471), .A1 (nx473), .A2 (nx475), .A3 (nx477)
           ) ;
    aoi22 ix472 (.Y (nx471), .A0 (x5[7]), .A1 (nx68), .B0 (x14[7]), .B1 (nx60)
          ) ;
    aoi22 ix474 (.Y (nx473), .A0 (x13[7]), .A1 (nx54), .B0 (x9[7]), .B1 (nx48)
          ) ;
    aoi22 ix476 (.Y (nx475), .A0 (x3[7]), .A1 (nx32), .B0 (x2[7]), .B1 (nx36)) ;
    aoi22 ix478 (.Y (nx477), .A0 (x8[7]), .A1 (nx10), .B0 (x10[7]), .B1 (nx18)
          ) ;
    buf02 ix483 (.Y (nx484), .A (nx78)) ;
    buf02 ix485 (.Y (nx486), .A (nx78)) ;
    inv02 ix491 (.Y (nx492), .A (nx261)) ;
    inv02 ix493 (.Y (nx495), .A (nx273)) ;
    inv02 ix496 (.Y (nx497), .A (nx295)) ;
    inv02 ix498 (.Y (nx499), .A (nx279)) ;
endmodule


module nbit_adder_12 ( a, b, cin, add_out ) ;

    input [11:0]a ;
    input [11:0]b ;
    input cin ;
    output [11:0]add_out ;

    wire temp_10, temp_9, temp_8, temp_7, temp_6, temp_5, temp_4, temp_3, temp_2, 
         temp_1, temp_0;
    wire [0:0] \$dummy ;




    bit_adder f0 (.a (a[0]), .b (b[0]), .cin (cin), .s (add_out[0]), .cout (
              temp_0)) ;
    bit_adder loop1_1_fx (.a (a[1]), .b (b[1]), .cin (temp_0), .s (add_out[1]), 
              .cout (temp_1)) ;
    bit_adder loop1_2_fx (.a (a[2]), .b (b[2]), .cin (temp_1), .s (add_out[2]), 
              .cout (temp_2)) ;
    bit_adder loop1_3_fx (.a (a[3]), .b (b[3]), .cin (temp_2), .s (add_out[3]), 
              .cout (temp_3)) ;
    bit_adder loop1_4_fx (.a (a[4]), .b (b[4]), .cin (temp_3), .s (add_out[4]), 
              .cout (temp_4)) ;
    bit_adder loop1_5_fx (.a (a[5]), .b (b[5]), .cin (temp_4), .s (add_out[5]), 
              .cout (temp_5)) ;
    bit_adder loop1_6_fx (.a (a[6]), .b (b[6]), .cin (temp_5), .s (add_out[6]), 
              .cout (temp_6)) ;
    bit_adder loop1_7_fx (.a (a[7]), .b (b[7]), .cin (temp_6), .s (add_out[7]), 
              .cout (temp_7)) ;
    bit_adder loop1_8_fx (.a (a[8]), .b (b[8]), .cin (temp_7), .s (add_out[8]), 
              .cout (temp_8)) ;
    bit_adder loop1_9_fx (.a (a[9]), .b (b[9]), .cin (temp_8), .s (add_out[9]), 
              .cout (temp_9)) ;
    bit_adder loop1_10_fx (.a (a[10]), .b (b[10]), .cin (temp_9), .s (
              add_out[10]), .cout (temp_10)) ;
    bit_adder loop1_11_fx (.a (a[11]), .b (b[11]), .cin (temp_10), .s (
              add_out[11]), .cout (\$dummy [0])) ;
endmodule


module DMACU ( clk, reset, start_DMA, Rows_Done, Row_Done, signals ) ;

    input clk ;
    input reset ;
    input start_DMA ;
    input Rows_Done ;
    input Row_Done ;
    output [5:0]signals ;

    wire state_4, state_1, nx4, nx12, nx28, nx40, nx62, nx74, nx224, nx226, 
         nx236, nx238, nx240, nx243;
    wire [5:0] \$dummy ;




    assign signals[2] = signals[5] ;
    or02 ix83 (.Y (signals[3]), .A0 (signals[4]), .A1 (state_4)) ;
    dff reg_state_2 (.Q (signals[4]), .QB (\$dummy [0]), .D (nx40), .CLK (clk)
        ) ;
    and03 ix41 (.Y (nx40), .A0 (state_1), .A1 (nx243), .A2 (start_DMA)) ;
    dff reg_state_1 (.Q (state_1), .QB (\$dummy [1]), .D (nx28), .CLK (clk)) ;
    nor02_2x ix29 (.Y (nx28), .A0 (reset), .A1 (nx224)) ;
    aoi21 ix225 (.Y (nx224), .A0 (nx226), .A1 (state_1), .B0 (signals[1])) ;
    inv01 ix227 (.Y (nx226), .A (start_DMA)) ;
    dff reg_state_0 (.Q (signals[1]), .QB (\$dummy [2]), .D (nx12), .CLK (clk)
        ) ;
    or02 ix13 (.Y (nx12), .A0 (signals[0]), .A1 (reset)) ;
    dff reg_state_5 (.Q (signals[0]), .QB (\$dummy [3]), .D (nx4), .CLK (clk)) ;
    and03 ix5 (.Y (nx4), .A0 (state_4), .A1 (nx243), .A2 (Rows_Done)) ;
    dff reg_state_4 (.Q (state_4), .QB (\$dummy [4]), .D (nx74), .CLK (clk)) ;
    and03 ix75 (.Y (nx74), .A0 (signals[5]), .A1 (nx243), .A2 (Row_Done)) ;
    dff reg_state_3 (.Q (signals[5]), .QB (\$dummy [5]), .D (nx62), .CLK (clk)
        ) ;
    nor02_2x ix63 (.Y (nx62), .A0 (reset), .A1 (nx236)) ;
    aoi221 ix237 (.Y (nx236), .A0 (nx238), .A1 (state_4), .B0 (nx240), .B1 (
           signals[5]), .C0 (signals[4])) ;
    inv01 ix239 (.Y (nx238), .A (Rows_Done)) ;
    inv01 ix241 (.Y (nx240), .A (Row_Done)) ;
    inv01 ix244 (.Y (nx243), .A (reset)) ;
endmodule


module \module  ( clk, rst, ack, start, move_done, nvm_address_in, cache_data_in, 
                  zero, one, cache_address_out, move, start_dma, done, direction, 
                  nvm_address_out, state_out ) ;

    input clk ;
    input rst ;
    input ack ;
    input start ;
    input move_done ;
    input [11:0]nvm_address_in ;
    input [7:0]cache_data_in ;
    input zero ;
    input one ;
    output [7:0]cache_address_out ;
    output move ;
    output start_dma ;
    output done ;
    output [0:0]direction ;
    output [11:0]nvm_address_out ;
    output [4:0]state_out ;

    wire pixel_value_17, pixel_value_16, pixel_value_15, pixel_value_14, 
         pixel_value_13, pixel_value_12, pixel_value_11, pixel_value_10, 
         pixel_value_9, pixel_value_8, pixel_value_7, pixel_value_6, 
         pixel_value_5, pixel_value_4, pixel_value_3, pixel_value_2, 
         pixel_value_1, pixel_value_0, sub_module_value_17, sub_module_value_16, 
         sub_module_value_15, sub_module_value_14, sub_module_value_13, 
         sub_module_value_12, sub_module_value_11, sub_module_value_10, 
         sub_module_value_9, sub_module_value_8, sub_module_value_7, 
         sub_module_value_6, sub_module_value_5, sub_module_value_4, 
         sub_module_value_3, sub_module_value_2, sub_module_value_1, 
         sub_module_value_0, bus_value_7, bus_value_6, bus_value_5, bus_value_4, 
         bus_value_3, bus_value_2, bus_value_1, bus_value_0, diff_value_17, 
         diff_value_16, diff_value_15, diff_value_14, diff_value_13, 
         diff_value_12, diff_value_11, diff_value_10, diff_value_9, diff_value_8, 
         diff_value_7, diff_value_6, diff_value_5, diff_value_4, diff_value_3, 
         diff_value_2, diff_value_1, diff_value_0, current_cont_value_17, 
         current_cont_value_16, current_cont_value_15, current_cont_value_14, 
         current_cont_value_13, current_cont_value_12, current_cont_value_11, 
         current_cont_value_10, current_cont_value_9, current_cont_value_8, 
         current_cont_value_7, current_cont_value_6, current_cont_value_5, 
         current_cont_value_4, current_cont_value_3, current_cont_value_2, 
         current_cont_value_1, current_cont_value_0, prev_cont_value_17, 
         prev_cont_value_16, prev_cont_value_15, prev_cont_value_14, 
         prev_cont_value_13, prev_cont_value_12, prev_cont_value_11, 
         prev_cont_value_10, prev_cont_value_9, prev_cont_value_8, 
         prev_cont_value_7, prev_cont_value_6, prev_cont_value_5, 
         prev_cont_value_4, prev_cont_value_3, prev_cont_value_2, 
         prev_cont_value_1, prev_cont_value_0, Addout_value_17, Addout_value_16, 
         Addout_value_15, Addout_value_14, Addout_value_13, Addout_value_12, 
         Addout_value_11, Addout_value_10, Addout_value_9, Addout_value_8, 
         Addout_value_7, Addout_value_6, Addout_value_5, Addout_value_4, 
         Addout_value_3, Addout_value_2, Addout_value_1, Addout_value_0, 
         add_module_value_17, add_module_value_16, add_module_value_15, 
         add_module_value_14, add_module_value_13, add_module_value_12, 
         add_module_value_11, add_module_value_10, add_module_value_9, 
         add_module_value_8, add_module_value_7, add_module_value_6, 
         add_module_value_5, add_module_value_4, add_module_value_3, 
         add_module_value_2, add_module_value_1, add_module_value_0, 
         prev_cont_bar_17, prev_cont_bar_16, prev_cont_bar_15, prev_cont_bar_14, 
         prev_cont_bar_13, prev_cont_bar_12, prev_cont_bar_11, prev_cont_bar_10, 
         prev_cont_bar_9, prev_cont_bar_8, prev_cont_bar_7, prev_cont_bar_6, 
         prev_cont_bar_5, prev_cont_bar_4, prev_cont_bar_3, prev_cont_bar_2, 
         prev_cont_bar_1, prev_cont_bar_0, comp_fake_value_16, address_value_7, 
         address_value_6, address_value_5, address_value_4, address_value_3, 
         address_value_2, address_value_1, address_value_0, plus_minus1_value_7, 
         plus_minus1_value_6, plus_minus1_value_5, plus_minus1_value_4, 
         plus_minus1_value_3, plus_minus1_value_2, plus_minus1_value_1, 
         plus_minus1_value_0, plus_minus16_value_7, plus_minus16_value_6, 
         plus_minus16_value_5, plus_minus16_value_4, plus_minus16_value_3, 
         plus_minus16_value_2, plus_minus16_value_1, plus_minus16_value_0, 
         finish, mux1_sel, direc_value_bar_0, mux2_sel_1, mux2_sel_0, inc_dec, 
         address_enable, current_cont_enable, pixel_enable, prev_cont_enable, 
         Addout_enable, diff_enable, failure_count_enable, regs_rst, lap_rst, 
         failure_count_value_0, nx12, nx26, nx818, nx820, nx822, nx824, nx826, 
         nx828, nx830, nx832, nx834, nx836, nx838, nx840, nx842, nx844;
    wire [17:0] \$dummy ;




    nbit_Register_18 pixel_reg (.Clk (clk), .rst (nx842), .enable (pixel_enable)
                     , .d ({zero,zero,zero,zero,zero,zero,zero,zero,zero,zero,
                     bus_value_7,bus_value_6,bus_value_5,bus_value_4,bus_value_3
                     ,bus_value_2,bus_value_1,bus_value_0}), .rst_value ({zero,
                     zero,zero,zero,zero,zero,zero,zero,zero,zero,zero,zero,zero
                     ,zero,zero,zero,zero,zero}), .q ({pixel_value_17,
                     pixel_value_16,pixel_value_15,pixel_value_14,pixel_value_13
                     ,pixel_value_12,pixel_value_11,pixel_value_10,pixel_value_9
                     ,pixel_value_8,pixel_value_7,pixel_value_6,pixel_value_5,
                     pixel_value_4,pixel_value_3,pixel_value_2,pixel_value_1,
                     pixel_value_0})) ;
    nbit_Register_18 diff_reg (.Clk (clk), .rst (nx842), .enable (diff_enable), 
                     .d ({sub_module_value_17,sub_module_value_16,
                     sub_module_value_15,sub_module_value_14,sub_module_value_13
                     ,sub_module_value_12,sub_module_value_11,
                     sub_module_value_10,sub_module_value_9,sub_module_value_8,
                     sub_module_value_7,sub_module_value_6,sub_module_value_5,
                     sub_module_value_4,sub_module_value_3,sub_module_value_2,
                     sub_module_value_1,sub_module_value_0}), .rst_value ({zero,
                     zero,zero,zero,zero,zero,zero,zero,zero,zero,zero,zero,zero
                     ,zero,zero,zero,zero,zero}), .q ({diff_value_17,
                     diff_value_16,diff_value_15,diff_value_14,diff_value_13,
                     diff_value_12,diff_value_11,diff_value_10,diff_value_9,
                     diff_value_8,diff_value_7,diff_value_6,diff_value_5,
                     diff_value_4,diff_value_3,diff_value_2,diff_value_1,
                     diff_value_0})) ;
    nbit_Register_18 Addout_reg (.Clk (clk), .rst (nx842), .enable (
                     Addout_enable), .d ({add_module_value_17,
                     add_module_value_16,add_module_value_15,add_module_value_14
                     ,add_module_value_13,add_module_value_12,
                     add_module_value_11,add_module_value_10,add_module_value_9,
                     add_module_value_8,add_module_value_7,add_module_value_6,
                     add_module_value_5,add_module_value_4,add_module_value_3,
                     add_module_value_2,add_module_value_1,add_module_value_0})
                     , .rst_value ({zero,zero,zero,zero,zero,zero,zero,zero,zero
                     ,zero,zero,zero,zero,zero,zero,zero,zero,zero}), .q ({
                     Addout_value_17,Addout_value_16,Addout_value_15,
                     Addout_value_14,Addout_value_13,Addout_value_12,
                     Addout_value_11,Addout_value_10,Addout_value_9,
                     Addout_value_8,Addout_value_7,Addout_value_6,Addout_value_5
                     ,Addout_value_4,Addout_value_3,Addout_value_2,
                     Addout_value_1,Addout_value_0})) ;
    nbit_Register_18 curr_cont_reg (.Clk (clk), .rst (lap_rst), .enable (
                     current_cont_enable), .d ({Addout_value_17,Addout_value_16,
                     Addout_value_15,Addout_value_14,Addout_value_13,
                     Addout_value_12,Addout_value_11,Addout_value_10,
                     Addout_value_9,Addout_value_8,Addout_value_7,Addout_value_6
                     ,Addout_value_5,Addout_value_4,Addout_value_3,
                     Addout_value_2,Addout_value_1,Addout_value_0}), .rst_value (
                     {zero,zero,zero,zero,zero,zero,zero,zero,zero,zero,zero,
                     zero,zero,zero,zero,zero,zero,zero}), .q ({
                     current_cont_value_17,current_cont_value_16,
                     current_cont_value_15,current_cont_value_14,
                     current_cont_value_13,current_cont_value_12,
                     current_cont_value_11,current_cont_value_10,
                     current_cont_value_9,current_cont_value_8,
                     current_cont_value_7,current_cont_value_6,
                     current_cont_value_5,current_cont_value_4,
                     current_cont_value_3,current_cont_value_2,
                     current_cont_value_1,current_cont_value_0})) ;
    nbit_Register_18 prev_cont_reg (.Clk (clk), .rst (nx842), .enable (
                     prev_cont_enable), .d ({current_cont_value_17,
                     current_cont_value_16,current_cont_value_15,
                     current_cont_value_14,current_cont_value_13,
                     current_cont_value_12,current_cont_value_11,
                     current_cont_value_10,current_cont_value_9,
                     current_cont_value_8,current_cont_value_7,
                     current_cont_value_6,current_cont_value_5,
                     current_cont_value_4,current_cont_value_3,
                     current_cont_value_2,current_cont_value_1,
                     current_cont_value_0}), .rst_value ({zero,zero,zero,zero,
                     zero,zero,zero,zero,zero,zero,zero,zero,zero,zero,zero,zero
                     ,zero,zero}), .q ({prev_cont_value_17,prev_cont_value_16,
                     prev_cont_value_15,prev_cont_value_14,prev_cont_value_13,
                     prev_cont_value_12,prev_cont_value_11,prev_cont_value_10,
                     prev_cont_value_9,prev_cont_value_8,prev_cont_value_7,
                     prev_cont_value_6,prev_cont_value_5,prev_cont_value_4,
                     prev_cont_value_3,prev_cont_value_2,prev_cont_value_1,
                     prev_cont_value_0})) ;
    nbit_Register_8 Address_reg (.Clk (clk), .rst (lap_rst), .enable (
                    address_enable), .d ({plus_minus1_value_7,
                    plus_minus1_value_6,plus_minus1_value_5,plus_minus1_value_4,
                    plus_minus1_value_3,plus_minus1_value_2,plus_minus1_value_1,
                    plus_minus1_value_0}), .rst_value ({zero,zero,zero,zero,zero
                    ,zero,zero,zero}), .q ({address_value_7,address_value_6,
                    address_value_5,address_value_4,address_value_3,
                    address_value_2,address_value_1,address_value_0})) ;
    nbit_Register_12 nvm_address_reg (.Clk (clk), .rst (nx842), .enable (
                     start_dma), .d ({nvm_address_in[11],nvm_address_in[10],
                     nvm_address_in[9],nvm_address_in[8],nvm_address_in[7],
                     nvm_address_in[6],nvm_address_in[5],nvm_address_in[4],
                     nvm_address_in[3],nvm_address_in[2],nvm_address_in[1],
                     nvm_address_in[0]}), .rst_value ({zero,zero,zero,zero,zero,
                     zero,zero,zero,zero,zero,zero,zero}), .q ({
                     nvm_address_out[11],nvm_address_out[10],nvm_address_out[9],
                     nvm_address_out[8],nvm_address_out[7],nvm_address_out[6],
                     nvm_address_out[5],nvm_address_out[4],nvm_address_out[3],
                     nvm_address_out[2],nvm_address_out[1],nvm_address_out[0]})
                     ) ;
    nbit_Register_1 direc_reg (.Clk (clk), .rst (nx844), .enable (
                    comp_fake_value_16), .d ({direc_value_bar_0}), .rst_value ({
                    zero}), .q ({direction[0]})) ;
    nbit_Register_1 fail_count_reg (.Clk (clk), .rst (nx844), .enable (
                    failure_count_enable), .d ({one}), .rst_value ({zero}), .q (
                    {failure_count_value_0})) ;
    nbit_mux3x1_8 mux2 (.input1 ({nx818,nx822,nx826,nx830,nx834,nx838,
                  address_value_1,address_value_0}), .input2 ({
                  plus_minus1_value_7,plus_minus1_value_6,plus_minus1_value_5,
                  plus_minus1_value_4,plus_minus1_value_3,plus_minus1_value_2,
                  plus_minus1_value_1,plus_minus1_value_0}), .input3 ({
                  plus_minus16_value_7,plus_minus16_value_6,plus_minus16_value_5
                  ,plus_minus16_value_4,plus_minus16_value_3,
                  plus_minus16_value_2,plus_minus16_value_1,plus_minus16_value_0
                  }), .s ({mux2_sel_1,mux2_sel_0}), .\output  ({
                  cache_address_out[7],cache_address_out[6],cache_address_out[5]
                  ,cache_address_out[4],cache_address_out[3],
                  cache_address_out[2],cache_address_out[1],cache_address_out[0]
                  })) ;
    nbit_mux2x1_8 mux1 (.input1 ({zero,zero,zero,zero,zero,zero,zero,zero}), .input2 (
                  {cache_data_in[7],cache_data_in[6],cache_data_in[5],
                  cache_data_in[4],cache_data_in[3],cache_data_in[2],
                  cache_data_in[1],cache_data_in[0]}), .s0 (mux1_sel), .\output  (
                  {bus_value_7,bus_value_6,bus_value_5,bus_value_4,bus_value_3,
                  bus_value_2,bus_value_1,bus_value_0})) ;
    selectData mux1_sel_block (.inc_dec (inc_dec), .s ({mux2_sel_1,mux2_sel_0})
               , .address ({nx818,nx822,nx826,nx830,nx834,nx838,address_value_1,
               address_value_0}), .func (mux1_sel)) ;
    sub submodule (.A ({pixel_value_17,pixel_value_16,pixel_value_15,
        pixel_value_14,pixel_value_13,pixel_value_12,pixel_value_11,
        pixel_value_10,pixel_value_9,pixel_value_8,pixel_value_7,pixel_value_6,
        pixel_value_5,pixel_value_4,pixel_value_3,pixel_value_2,pixel_value_1,
        pixel_value_0}), .B ({zero,zero,zero,zero,zero,zero,zero,zero,zero,zero,
        bus_value_7,bus_value_6,bus_value_5,bus_value_4,bus_value_3,bus_value_2,
        bus_value_1,bus_value_0}), .zero (zero), .one (one), .sub_value ({
        sub_module_value_17,sub_module_value_16,sub_module_value_15,
        sub_module_value_14,sub_module_value_13,sub_module_value_12,
        sub_module_value_11,sub_module_value_10,sub_module_value_9,
        sub_module_value_8,sub_module_value_7,sub_module_value_6,
        sub_module_value_5,sub_module_value_4,sub_module_value_3,
        sub_module_value_2,sub_module_value_1,sub_module_value_0})) ;
    nbit_adder_18 addmodule (.a ({current_cont_value_17,current_cont_value_16,
                  current_cont_value_15,current_cont_value_14,
                  current_cont_value_13,current_cont_value_12,
                  current_cont_value_11,current_cont_value_10,
                  current_cont_value_9,current_cont_value_8,current_cont_value_7
                  ,current_cont_value_6,current_cont_value_5,
                  current_cont_value_4,current_cont_value_3,current_cont_value_2
                  ,current_cont_value_1,current_cont_value_0}), .b ({
                  diff_value_17,diff_value_16,diff_value_15,diff_value_14,
                  diff_value_13,diff_value_12,diff_value_11,diff_value_10,
                  diff_value_9,diff_value_8,diff_value_7,diff_value_6,
                  diff_value_5,diff_value_4,diff_value_3,diff_value_2,
                  diff_value_1,diff_value_0}), .cin (zero), .add_out ({
                  add_module_value_17,add_module_value_16,add_module_value_15,
                  add_module_value_14,add_module_value_13,add_module_value_12,
                  add_module_value_11,add_module_value_10,add_module_value_9,
                  add_module_value_8,add_module_value_7,add_module_value_6,
                  add_module_value_5,add_module_value_4,add_module_value_3,
                  add_module_value_2,add_module_value_1,add_module_value_0})) ;
    nbit_adder_18 compmodule (.a ({current_cont_value_17,current_cont_value_16,
                  current_cont_value_15,current_cont_value_14,
                  current_cont_value_13,current_cont_value_12,
                  current_cont_value_11,current_cont_value_10,
                  current_cont_value_9,current_cont_value_8,current_cont_value_7
                  ,current_cont_value_6,current_cont_value_5,
                  current_cont_value_4,current_cont_value_3,current_cont_value_2
                  ,current_cont_value_1,current_cont_value_0}), .b ({
                  prev_cont_bar_17,prev_cont_bar_16,prev_cont_bar_15,
                  prev_cont_bar_14,prev_cont_bar_13,prev_cont_bar_12,
                  prev_cont_bar_11,prev_cont_bar_10,prev_cont_bar_9,
                  prev_cont_bar_8,prev_cont_bar_7,prev_cont_bar_6,
                  prev_cont_bar_5,prev_cont_bar_4,prev_cont_bar_3,
                  prev_cont_bar_2,prev_cont_bar_1,prev_cont_bar_0}), .cin (one)
                  , .add_out ({\$dummy [0],comp_fake_value_16,\$dummy [1],
                  \$dummy [2],\$dummy [3],\$dummy [4],\$dummy [5],\$dummy [6],
                  \$dummy [7],\$dummy [8],\$dummy [9],\$dummy [10],\$dummy [11],
                  \$dummy [12],\$dummy [13],\$dummy [14],\$dummy [15],
                  \$dummy [16]})) ;
    inc_dec_module plusMinus1 (.A ({nx818,nx822,nx826,nx830,nx834,nx838,
                   address_value_1,address_value_0}), .amount ({zero,zero,zero,
                   zero,zero,zero,zero,one}), .inc_dec (inc_dec), .\output  ({
                   plus_minus1_value_7,plus_minus1_value_6,plus_minus1_value_5,
                   plus_minus1_value_4,plus_minus1_value_3,plus_minus1_value_2,
                   plus_minus1_value_1,plus_minus1_value_0})) ;
    inc_dec_module plusMinus16 (.A ({nx818,nx822,nx826,nx830,nx834,nx838,
                   address_value_1,address_value_0}), .amount ({zero,zero,zero,
                   one,zero,zero,zero,zero}), .inc_dec (inc_dec), .\output  ({
                   plus_minus16_value_7,plus_minus16_value_6,
                   plus_minus16_value_5,plus_minus16_value_4,
                   plus_minus16_value_3,plus_minus16_value_2,
                   plus_minus16_value_1,plus_minus16_value_0})) ;
    module_CU modCU (.\input  ({failure_count_value_0,comp_fake_value_16,
              move_done,start,ack,finish}), .signals ({lap_rst,regs_rst,
              mux2_sel_1,mux2_sel_0,inc_dec,address_enable,current_cont_enable,
              pixel_enable,prev_cont_enable,Addout_enable,diff_enable,start_dma,
              move,\$dummy [17],done,failure_count_enable}), .state_out ({
              state_out[4],state_out[3],state_out[2],state_out[1],state_out[0]})
              , .clk (clk), .rst_sig (rst)) ;
    inv01 ix773 (.Y (direc_value_bar_0), .A (direction[0])) ;
    and02 ix29 (.Y (finish), .A0 (nx12), .A1 (nx26)) ;
    nor04 ix13 (.Y (nx12), .A0 (address_value_0), .A1 (address_value_1), .A2 (
          nx840), .A3 (nx836)) ;
    nor04 ix27 (.Y (nx26), .A0 (nx832), .A1 (nx828), .A2 (nx824), .A3 (nx820)) ;
    inv01 ix778 (.Y (prev_cont_bar_0), .A (prev_cont_value_0)) ;
    inv01 ix780 (.Y (prev_cont_bar_1), .A (prev_cont_value_1)) ;
    inv01 ix782 (.Y (prev_cont_bar_2), .A (prev_cont_value_2)) ;
    inv01 ix784 (.Y (prev_cont_bar_3), .A (prev_cont_value_3)) ;
    inv01 ix786 (.Y (prev_cont_bar_4), .A (prev_cont_value_4)) ;
    inv01 ix788 (.Y (prev_cont_bar_5), .A (prev_cont_value_5)) ;
    inv01 ix790 (.Y (prev_cont_bar_6), .A (prev_cont_value_6)) ;
    inv01 ix792 (.Y (prev_cont_bar_7), .A (prev_cont_value_7)) ;
    inv01 ix794 (.Y (prev_cont_bar_8), .A (prev_cont_value_8)) ;
    inv01 ix796 (.Y (prev_cont_bar_9), .A (prev_cont_value_9)) ;
    inv01 ix798 (.Y (prev_cont_bar_10), .A (prev_cont_value_10)) ;
    inv01 ix800 (.Y (prev_cont_bar_11), .A (prev_cont_value_11)) ;
    inv01 ix802 (.Y (prev_cont_bar_12), .A (prev_cont_value_12)) ;
    inv01 ix804 (.Y (prev_cont_bar_13), .A (prev_cont_value_13)) ;
    inv01 ix806 (.Y (prev_cont_bar_14), .A (prev_cont_value_14)) ;
    inv01 ix808 (.Y (prev_cont_bar_15), .A (prev_cont_value_15)) ;
    inv01 ix810 (.Y (prev_cont_bar_16), .A (prev_cont_value_16)) ;
    inv01 ix812 (.Y (prev_cont_bar_17), .A (prev_cont_value_17)) ;
    buf02 ix817 (.Y (nx818), .A (address_value_7)) ;
    buf02 ix819 (.Y (nx820), .A (address_value_7)) ;
    buf02 ix821 (.Y (nx822), .A (address_value_6)) ;
    buf02 ix823 (.Y (nx824), .A (address_value_6)) ;
    buf02 ix825 (.Y (nx826), .A (address_value_5)) ;
    buf02 ix827 (.Y (nx828), .A (address_value_5)) ;
    buf02 ix829 (.Y (nx830), .A (address_value_4)) ;
    buf02 ix831 (.Y (nx832), .A (address_value_4)) ;
    buf02 ix833 (.Y (nx834), .A (address_value_3)) ;
    buf02 ix835 (.Y (nx836), .A (address_value_3)) ;
    buf02 ix837 (.Y (nx838), .A (address_value_2)) ;
    buf02 ix839 (.Y (nx840), .A (address_value_2)) ;
    buf02 ix841 (.Y (nx842), .A (regs_rst)) ;
    buf02 ix843 (.Y (nx844), .A (regs_rst)) ;
endmodule


module module_CU ( \input , signals, state_out, clk, rst_sig ) ;

    input [5:0]\input  ;
    output [15:0]signals ;
    output [4:0]state_out ;
    input clk ;
    input rst_sig ;

    wire current_state_13, nx705, current_state_10, current_state_9, 
         current_state_8, current_state_7, current_state_6, current_state_4, 
         current_state_14, nx20, nx24, current_state_1, nx56, nx80, 
         current_state_12, nx108, nx188, nx226, nx294, nx710, nx722, nx732, 
         nx742, nx752, nx762, nx772, nx780, nx792, nx802, nx812, nx822, nx832, 
         nx842, nx852, nx862, nx872, nx880, nx893, nx902, nx906, nx910, nx913, 
         nx915, nx922, nx928, nx939, nx942, nx946, nx948, nx952, nx954, nx959, 
         nx964, nx968, nx970, nx973, nx977, nx980, nx984, nx986, nx988, nx993, 
         nx995, nx998, nx1000, nx1004, nx1010, nx1012, nx1016, nx1018, nx1021, 
         nx1023, nx1025, nx1027, nx1036, nx1038, nx1040, nx1042, nx1044, nx1052, 
         nx1054, nx1056, nx1058, nx1060, nx1062;
    wire [7:0] \$dummy ;




    assign signals[2] = signals[4] ;
    nand03 ix283 (.Y (state_out[3]), .A0 (nx893), .A1 (nx977), .A2 (nx1004)) ;
    dff reg_current_state_11 (.Q (signals[10]), .QB (\$dummy [0]), .D (nx872), .CLK (
        clk)) ;
    dff reg_current_state_10 (.Q (current_state_10), .QB (nx902), .D (nx862), .CLK (
        clk)) ;
    oai21 ix863 (.Y (nx862), .A0 (nx902), .A1 (nx1040), .B0 (nx1000)) ;
    nand04 ix235 (.Y (nx705), .A0 (nx906), .A1 (nx928), .A2 (nx954), .A3 (nx988)
           ) ;
    nor04 ix907 (.Y (nx906), .A0 (current_state_13), .A1 (current_state_14), .A2 (
          rst_sig), .A3 (nx226)) ;
    dff reg_current_state_13 (.Q (current_state_13), .QB (nx910), .D (nx880), .CLK (
        clk)) ;
    dff reg_current_state_14 (.Q (current_state_14), .QB (nx913), .D (nx710), .CLK (
        clk)) ;
    nand03 ix227 (.Y (nx226), .A0 (nx915), .A1 (nx922), .A2 (nx998)) ;
    nand03 ix916 (.Y (nx915), .A0 (signals[3]), .A1 (nx1042), .A2 (\input [3])
           ) ;
    dff reg_current_state_15 (.Q (signals[3]), .QB (\$dummy [1]), .D (nx722), .CLK (
        clk)) ;
    nor02ii ix25 (.Y (nx24), .A0 (rst_sig), .A1 (nx20)) ;
    oai22 ix21 (.Y (nx20), .A0 (\input [5]), .A1 (nx913), .B0 (\input [4]), .B1 (
          nx910)) ;
    nor02_2x ix923 (.Y (nx922), .A0 (signals[7]), .A1 (signals[1])) ;
    dff reg_current_state_16 (.Q (signals[7]), .QB (\$dummy [2]), .D (nx732), .CLK (
        clk)) ;
    ao32 ix733 (.Y (nx732), .A0 (signals[3]), .A1 (nx1042), .A2 (\input [3]), .B0 (
         signals[7]), .B1 (nx1058)) ;
    aoi21 ix929 (.Y (nx928), .A0 (nx1042), .A1 (signals[14]), .B0 (signals[5])
          ) ;
    dff reg_current_state_0 (.Q (signals[14]), .QB (\$dummy [3]), .D (nx752), .CLK (
        clk)) ;
    or02 ix57 (.Y (nx56), .A0 (signals[1]), .A1 (rst_sig)) ;
    dff reg_current_state_17 (.Q (signals[1]), .QB (\$dummy [4]), .D (nx742), .CLK (
        clk)) ;
    ao32 ix743 (.Y (nx742), .A0 (current_state_14), .A1 (nx1042), .A2 (
         \input [5]), .B0 (signals[1]), .B1 (nx1058)) ;
    or02 ix215 (.Y (signals[5]), .A0 (signals[13]), .A1 (signals[12])) ;
    dff reg_current_state_6 (.Q (current_state_6), .QB (nx939), .D (nx822), .CLK (
        clk)) ;
    oai21 ix823 (.Y (nx822), .A0 (nx939), .A1 (nx1036), .B0 (nx942)) ;
    oai21 ix813 (.Y (nx812), .A0 (nx946), .A1 (nx1036), .B0 (nx948)) ;
    dff reg_current_state_5 (.Q (\$dummy [5]), .QB (nx946), .D (nx812), .CLK (
        clk)) ;
    oai21 ix803 (.Y (nx802), .A0 (nx952), .A1 (nx1036), .B0 (nx954)) ;
    dff reg_current_state_4 (.Q (current_state_4), .QB (nx952), .D (nx802), .CLK (
        clk)) ;
    nand02 ix955 (.Y (nx954), .A0 (nx1044), .A1 (signals[8])) ;
    dff reg_current_state_3 (.Q (signals[8]), .QB (\$dummy [6]), .D (nx792), .CLK (
        clk)) ;
    nor02_2x ix109 (.Y (nx108), .A0 (rst_sig), .A1 (nx959)) ;
    aoi22 ix960 (.Y (nx959), .A0 (\input [1]), .A1 (signals[4]), .B0 (nx973), .B1 (
          current_state_12)) ;
    dff reg_current_state_2 (.Q (signals[4]), .QB (\$dummy [7]), .D (nx772), .CLK (
        clk)) ;
    nor02_2x ix81 (.Y (nx80), .A0 (rst_sig), .A1 (nx964)) ;
    aoi21 ix965 (.Y (nx964), .A0 (\input [2]), .A1 (current_state_1), .B0 (
          signals[7])) ;
    oai21 ix763 (.Y (nx762), .A0 (nx968), .A1 (nx1036), .B0 (nx970)) ;
    dff reg_current_state_1 (.Q (current_state_1), .QB (nx968), .D (nx762), .CLK (
        clk)) ;
    nand02 ix971 (.Y (nx970), .A0 (nx1044), .A1 (signals[14])) ;
    inv01 ix974 (.Y (nx973), .A (\input [0])) ;
    dff reg_current_state_8 (.Q (current_state_8), .QB (nx977), .D (nx842), .CLK (
        clk)) ;
    oai21 ix843 (.Y (nx842), .A0 (nx977), .A1 (nx1038), .B0 (nx980)) ;
    oai21 ix833 (.Y (nx832), .A0 (nx984), .A1 (nx1038), .B0 (nx986)) ;
    dff reg_current_state_7 (.Q (current_state_7), .QB (nx984), .D (nx832), .CLK (
        clk)) ;
    aoi221 ix989 (.Y (nx988), .A0 (\input [1]), .A1 (signals[4]), .B0 (
           \input [2]), .B1 (current_state_1), .C0 (signals[6])) ;
    oai21 ix853 (.Y (nx852), .A0 (nx993), .A1 (nx1040), .B0 (nx995)) ;
    dff reg_current_state_9 (.Q (current_state_9), .QB (nx993), .D (nx852), .CLK (
        clk)) ;
    dff reg_current_state_12 (.Q (current_state_12), .QB (nx998), .D (nx780), .CLK (
        clk)) ;
    nor03_2x ix1005 (.Y (nx1004), .A0 (current_state_10), .A1 (signals[10]), .A2 (
             current_state_9)) ;
    or02 ix311 (.Y (signals[15]), .A0 (signals[14]), .A1 (signals[7])) ;
    nand02 ix257 (.Y (state_out[0]), .A0 (nx1010), .A1 (nx1012)) ;
    nor03_2x ix1011 (.Y (nx1010), .A0 (current_state_1), .A1 (signals[8]), .A2 (
             signals[6])) ;
    nor03_2x ix1013 (.Y (nx1012), .A0 (signals[3]), .A1 (signals[7]), .A2 (
             current_state_13)) ;
    nand04 ix303 (.Y (state_out[1]), .A0 (nx294), .A1 (nx1023), .A2 (nx1025), .A3 (
           nx1027)) ;
    nand04 ix295 (.Y (nx294), .A0 (nx1016), .A1 (nx922), .A2 (nx1018), .A3 (
           nx1021)) ;
    nor04 ix1022 (.Y (nx1021), .A0 (signals[14]), .A1 (current_state_1), .A2 (
          signals[4]), .A3 (signals[8])) ;
    nor04 ix1028 (.Y (nx1027), .A0 (signals[4]), .A1 (signals[8]), .A2 (
          current_state_7), .A3 (signals[10])) ;
    nand02 ix313 (.Y (state_out[2]), .A0 (nx893), .A1 (nx1016)) ;
    nand02 ix317 (.Y (state_out[4]), .A0 (nx294), .A1 (nx922)) ;
    inv01 ix1019 (.Y (nx1018), .A (state_out[3])) ;
    inv01 ix265 (.Y (signals[0]), .A (nx1023)) ;
    inv01 ix213 (.Y (signals[13]), .A (nx1025)) ;
    inv02 ix1035 (.Y (nx1036), .A (nx1058)) ;
    inv02 ix1037 (.Y (nx1038), .A (nx1058)) ;
    inv02 ix1039 (.Y (nx1040), .A (nx1058)) ;
    inv02 ix1041 (.Y (nx1042), .A (rst_sig)) ;
    inv02 ix1043 (.Y (nx1044), .A (rst_sig)) ;
    and03 ix894 (.Y (nx893), .A0 (nx998), .A1 (nx910), .A2 (nx1023)) ;
    nor03_2x ix781 (.Y (nx780), .A0 (rst_sig), .A1 (nx1052), .A2 (nx1058)) ;
    inv01 ix1051 (.Y (nx1052), .A (signals[10])) ;
    mux21_ni ix873 (.Y (nx872), .A0 (nx188), .A1 (signals[10]), .S0 (nx1058)) ;
    nor02ii ix189 (.Y (nx188), .A0 (rst_sig), .A1 (current_state_10)) ;
    nor03_2x ix881 (.Y (nx880), .A0 (nx998), .A1 (rst_sig), .A2 (nx973)) ;
    nor03_2x ix711 (.Y (nx710), .A0 (nx910), .A1 (rst_sig), .A2 (nx1054)) ;
    inv01 ix1053 (.Y (nx1054), .A (\input [4])) ;
    mux21_ni ix723 (.Y (nx722), .A0 (nx24), .A1 (signals[3]), .S0 (nx1060)) ;
    mux21_ni ix753 (.Y (nx752), .A0 (nx56), .A1 (signals[14]), .S0 (nx1060)) ;
    or03 ix943 (.Y (nx942), .A0 (rst_sig), .A1 (nx946), .A2 (nx1060)) ;
    or03 ix949 (.Y (nx948), .A0 (rst_sig), .A1 (nx952), .A2 (nx1060)) ;
    mux21_ni ix793 (.Y (nx792), .A0 (nx108), .A1 (signals[8]), .S0 (nx1060)) ;
    mux21_ni ix773 (.Y (nx772), .A0 (nx80), .A1 (signals[4]), .S0 (nx1060)) ;
    or02 ix211 (.Y (signals[12]), .A0 (current_state_4), .A1 (current_state_8)
         ) ;
    or03 ix981 (.Y (nx980), .A0 (rst_sig), .A1 (nx984), .A2 (nx1060)) ;
    or03 ix987 (.Y (nx986), .A0 (rst_sig), .A1 (nx939), .A2 (nx1062)) ;
    nand04 ix201 (.Y (signals[6]), .A0 (nx946), .A1 (nx984), .A2 (nx993), .A3 (
           nx1052)) ;
    or03 ix996 (.Y (nx995), .A0 (rst_sig), .A1 (nx977), .A2 (nx1062)) ;
    or03 ix1001 (.Y (nx1000), .A0 (rst_sig), .A1 (nx993), .A2 (nx1062)) ;
    nand03 ix309 (.Y (signals[9]), .A0 (nx902), .A1 (nx998), .A2 (nx1056)) ;
    inv01 ix1055 (.Y (nx1056), .A (signals[11])) ;
    or02 ix305 (.Y (signals[11]), .A0 (current_state_6), .A1 (current_state_8)
         ) ;
    and04 ix1017 (.Y (nx1016), .A0 (nx952), .A1 (nx946), .A2 (nx939), .A3 (nx984
          )) ;
    nor02ii ix1024 (.Y (nx1023), .A0 (signals[3]), .A1 (nx913)) ;
    and02 ix1026 (.Y (nx1025), .A0 (nx939), .A1 (nx902)) ;
    inv02 ix1057 (.Y (nx1058), .A (nx705)) ;
    inv02 ix1059 (.Y (nx1060), .A (nx705)) ;
    inv02 ix1061 (.Y (nx1062), .A (nx705)) ;
endmodule


module inc_dec_module ( A, amount, inc_dec, \output  ) ;

    input [7:0]A ;
    input [7:0]amount ;
    input inc_dec ;
    output [7:0]\output  ;

    wire amount_to_adder_7, amount_to_adder_6, amount_to_adder_5, 
         amount_to_adder_4, amount_to_adder_3, amount_to_adder_2, 
         amount_to_adder_1, amount_to_adder_0, nx197, nx199, nx201;



    nbit_adder_8 u (.a ({A[7],A[6],A[5],A[4],A[3],A[2],A[1],A[0]}), .b ({
                 amount_to_adder_7,amount_to_adder_6,amount_to_adder_5,
                 amount_to_adder_4,amount_to_adder_3,amount_to_adder_2,
                 amount_to_adder_1,amount_to_adder_0}), .cin (nx199), .add_out (
                 {\output [7],\output [6],\output [5],\output [4],\output [3],
                 \output [2],\output [1],\output [0]})) ;
    xor2 ix1 (.Y (amount_to_adder_0), .A0 (amount[0]), .A1 (nx199)) ;
    xor2 ix3 (.Y (amount_to_adder_1), .A0 (amount[1]), .A1 (nx199)) ;
    xor2 ix5 (.Y (amount_to_adder_2), .A0 (amount[2]), .A1 (nx199)) ;
    xor2 ix7 (.Y (amount_to_adder_3), .A0 (amount[3]), .A1 (nx199)) ;
    xor2 ix9 (.Y (amount_to_adder_4), .A0 (amount[4]), .A1 (nx201)) ;
    xor2 ix11 (.Y (amount_to_adder_5), .A0 (amount[5]), .A1 (nx201)) ;
    xor2 ix13 (.Y (amount_to_adder_6), .A0 (amount[6]), .A1 (nx201)) ;
    xor2 ix15 (.Y (amount_to_adder_7), .A0 (amount[7]), .A1 (nx201)) ;
    inv01 ix196 (.Y (nx197), .A (inc_dec)) ;
    inv02 ix198 (.Y (nx199), .A (nx197)) ;
    inv02 ix200 (.Y (nx201), .A (nx197)) ;
endmodule


module nbit_adder_8 ( a, b, cin, add_out ) ;

    input [7:0]a ;
    input [7:0]b ;
    input cin ;
    output [7:0]add_out ;

    wire temp_6, temp_5, temp_4, temp_3, temp_2, temp_1, temp_0;
    wire [0:0] \$dummy ;




    bit_adder f0 (.a (a[0]), .b (b[0]), .cin (cin), .s (add_out[0]), .cout (
              temp_0)) ;
    bit_adder loop1_1_fx (.a (a[1]), .b (b[1]), .cin (temp_0), .s (add_out[1]), 
              .cout (temp_1)) ;
    bit_adder loop1_2_fx (.a (a[2]), .b (b[2]), .cin (temp_1), .s (add_out[2]), 
              .cout (temp_2)) ;
    bit_adder loop1_3_fx (.a (a[3]), .b (b[3]), .cin (temp_2), .s (add_out[3]), 
              .cout (temp_3)) ;
    bit_adder loop1_4_fx (.a (a[4]), .b (b[4]), .cin (temp_3), .s (add_out[4]), 
              .cout (temp_4)) ;
    bit_adder loop1_5_fx (.a (a[5]), .b (b[5]), .cin (temp_4), .s (add_out[5]), 
              .cout (temp_5)) ;
    bit_adder loop1_6_fx (.a (a[6]), .b (b[6]), .cin (temp_5), .s (add_out[6]), 
              .cout (temp_6)) ;
    bit_adder loop1_7_fx (.a (a[7]), .b (b[7]), .cin (temp_6), .s (add_out[7]), 
              .cout (\$dummy [0])) ;
endmodule


module sub ( A, B, zero, one, sub_value ) ;

    input [17:0]A ;
    input [17:0]B ;
    input zero ;
    input one ;
    output [17:0]sub_value ;

    wire B_bar_17, B_bar_16, B_bar_15, B_bar_14, B_bar_13, B_bar_12, B_bar_11, 
         B_bar_10, B_bar_9, B_bar_8, B_bar_7, B_bar_6, B_bar_5, B_bar_4, B_bar_3, 
         B_bar_2, B_bar_1, B_bar_0, Adder1_value_17, Adder1_value_16, 
         Adder1_value_15, Adder1_value_14, Adder1_value_13, Adder1_value_12, 
         Adder1_value_11, Adder1_value_10, Adder1_value_9, Adder1_value_8, 
         Adder1_value_7, Adder1_value_6, Adder1_value_5, Adder1_value_4, 
         Adder1_value_3, Adder1_value_2, Adder1_value_1, Adder1_value_0, 
         Adder2_value_17, Adder2_value_16, Adder2_value_15, Adder2_value_14, 
         Adder2_value_13, Adder2_value_12, Adder2_value_11, Adder2_value_10, 
         Adder2_value_9, Adder2_value_8, Adder2_value_7, Adder2_value_6, 
         Adder2_value_5, Adder2_value_4, Adder2_value_3, Adder2_value_2, 
         Adder2_value_1, Adder2_value_0, Adder1_value_bar_17, 
         Adder1_value_bar_15, Adder1_value_bar_14, Adder1_value_bar_13, 
         Adder1_value_bar_12, Adder1_value_bar_11, Adder1_value_bar_10, 
         Adder1_value_bar_9, Adder1_value_bar_8, Adder1_value_bar_7, 
         Adder1_value_bar_6, Adder1_value_bar_5, Adder1_value_bar_4, 
         Adder1_value_bar_3, Adder1_value_bar_2, Adder1_value_bar_1, 
         Adder1_value_bar_0, nx452, nx454, nx456;



    nbit_adder_18 Adder1_sub (.a ({A[17],A[16],A[15],A[14],A[13],A[12],A[11],
                  A[10],A[9],A[8],A[7],A[6],A[5],A[4],A[3],A[2],A[1],A[0]}), .b (
                  {B_bar_17,B_bar_16,B_bar_15,B_bar_14,B_bar_13,B_bar_12,
                  B_bar_11,B_bar_10,B_bar_9,B_bar_8,B_bar_7,B_bar_6,B_bar_5,
                  B_bar_4,B_bar_3,B_bar_2,B_bar_1,B_bar_0}), .cin (one), .add_out (
                  {Adder1_value_17,Adder1_value_16,Adder1_value_15,
                  Adder1_value_14,Adder1_value_13,Adder1_value_12,
                  Adder1_value_11,Adder1_value_10,Adder1_value_9,Adder1_value_8,
                  Adder1_value_7,Adder1_value_6,Adder1_value_5,Adder1_value_4,
                  Adder1_value_3,Adder1_value_2,Adder1_value_1,Adder1_value_0})
                  ) ;
    nbit_adder_18 Adder2_sub (.a ({Adder1_value_bar_17,nx452,Adder1_value_bar_15
                  ,Adder1_value_bar_14,Adder1_value_bar_13,Adder1_value_bar_12,
                  Adder1_value_bar_11,Adder1_value_bar_10,Adder1_value_bar_9,
                  Adder1_value_bar_8,Adder1_value_bar_7,Adder1_value_bar_6,
                  Adder1_value_bar_5,Adder1_value_bar_4,Adder1_value_bar_3,
                  Adder1_value_bar_2,Adder1_value_bar_1,Adder1_value_bar_0}), .b (
                  {zero,zero,zero,zero,zero,zero,zero,zero,zero,zero,zero,zero,
                  zero,zero,zero,zero,zero,zero}), .cin (one), .add_out ({
                  Adder2_value_17,Adder2_value_16,Adder2_value_15,
                  Adder2_value_14,Adder2_value_13,Adder2_value_12,
                  Adder2_value_11,Adder2_value_10,Adder2_value_9,Adder2_value_8,
                  Adder2_value_7,Adder2_value_6,Adder2_value_5,Adder2_value_4,
                  Adder2_value_3,Adder2_value_2,Adder2_value_1,Adder2_value_0})
                  ) ;
    inv01 ix348 (.Y (Adder1_value_bar_0), .A (Adder1_value_0)) ;
    inv01 ix350 (.Y (Adder1_value_bar_1), .A (Adder1_value_1)) ;
    inv01 ix352 (.Y (Adder1_value_bar_2), .A (Adder1_value_2)) ;
    inv01 ix354 (.Y (Adder1_value_bar_3), .A (Adder1_value_3)) ;
    inv01 ix356 (.Y (Adder1_value_bar_4), .A (Adder1_value_4)) ;
    inv01 ix358 (.Y (Adder1_value_bar_5), .A (Adder1_value_5)) ;
    inv01 ix360 (.Y (Adder1_value_bar_6), .A (Adder1_value_6)) ;
    inv01 ix362 (.Y (Adder1_value_bar_7), .A (Adder1_value_7)) ;
    inv01 ix364 (.Y (Adder1_value_bar_8), .A (Adder1_value_8)) ;
    inv01 ix366 (.Y (Adder1_value_bar_9), .A (Adder1_value_9)) ;
    inv01 ix368 (.Y (Adder1_value_bar_10), .A (Adder1_value_10)) ;
    inv01 ix370 (.Y (Adder1_value_bar_11), .A (Adder1_value_11)) ;
    inv01 ix372 (.Y (Adder1_value_bar_12), .A (Adder1_value_12)) ;
    inv01 ix374 (.Y (Adder1_value_bar_13), .A (Adder1_value_13)) ;
    inv01 ix376 (.Y (Adder1_value_bar_14), .A (Adder1_value_14)) ;
    inv01 ix378 (.Y (Adder1_value_bar_15), .A (Adder1_value_15)) ;
    inv01 ix382 (.Y (Adder1_value_bar_17), .A (Adder1_value_17)) ;
    inv01 ix402 (.Y (B_bar_0), .A (B[0])) ;
    inv01 ix404 (.Y (B_bar_1), .A (B[1])) ;
    inv01 ix406 (.Y (B_bar_2), .A (B[2])) ;
    inv01 ix408 (.Y (B_bar_3), .A (B[3])) ;
    inv01 ix410 (.Y (B_bar_4), .A (B[4])) ;
    inv01 ix412 (.Y (B_bar_5), .A (B[5])) ;
    inv01 ix414 (.Y (B_bar_6), .A (B[6])) ;
    inv01 ix416 (.Y (B_bar_7), .A (B[7])) ;
    inv01 ix418 (.Y (B_bar_8), .A (B[8])) ;
    inv01 ix420 (.Y (B_bar_9), .A (B[9])) ;
    inv01 ix422 (.Y (B_bar_10), .A (B[10])) ;
    inv01 ix424 (.Y (B_bar_11), .A (B[11])) ;
    inv01 ix426 (.Y (B_bar_12), .A (B[12])) ;
    inv01 ix428 (.Y (B_bar_13), .A (B[13])) ;
    inv01 ix430 (.Y (B_bar_14), .A (B[14])) ;
    inv01 ix432 (.Y (B_bar_15), .A (B[15])) ;
    inv01 ix434 (.Y (B_bar_16), .A (B[16])) ;
    inv01 ix436 (.Y (B_bar_17), .A (B[17])) ;
    mux21_ni ix9 (.Y (sub_value[0]), .A0 (Adder2_value_0), .A1 (Adder1_value_0)
             , .S0 (nx452)) ;
    mux21_ni ix17 (.Y (sub_value[1]), .A0 (Adder2_value_1), .A1 (Adder1_value_1)
             , .S0 (nx452)) ;
    mux21_ni ix25 (.Y (sub_value[2]), .A0 (Adder2_value_2), .A1 (Adder1_value_2)
             , .S0 (nx452)) ;
    mux21_ni ix33 (.Y (sub_value[3]), .A0 (Adder2_value_3), .A1 (Adder1_value_3)
             , .S0 (nx452)) ;
    mux21_ni ix41 (.Y (sub_value[4]), .A0 (Adder2_value_4), .A1 (Adder1_value_4)
             , .S0 (nx452)) ;
    mux21_ni ix49 (.Y (sub_value[5]), .A0 (Adder2_value_5), .A1 (Adder1_value_5)
             , .S0 (nx454)) ;
    mux21_ni ix57 (.Y (sub_value[6]), .A0 (Adder2_value_6), .A1 (Adder1_value_6)
             , .S0 (nx454)) ;
    mux21_ni ix65 (.Y (sub_value[7]), .A0 (Adder2_value_7), .A1 (Adder1_value_7)
             , .S0 (nx454)) ;
    mux21_ni ix73 (.Y (sub_value[8]), .A0 (Adder2_value_8), .A1 (Adder1_value_8)
             , .S0 (nx454)) ;
    mux21_ni ix81 (.Y (sub_value[9]), .A0 (Adder2_value_9), .A1 (Adder1_value_9)
             , .S0 (nx454)) ;
    mux21_ni ix89 (.Y (sub_value[10]), .A0 (Adder2_value_10), .A1 (
             Adder1_value_10), .S0 (nx454)) ;
    mux21_ni ix97 (.Y (sub_value[11]), .A0 (Adder2_value_11), .A1 (
             Adder1_value_11), .S0 (nx454)) ;
    mux21_ni ix105 (.Y (sub_value[12]), .A0 (Adder2_value_12), .A1 (
             Adder1_value_12), .S0 (nx456)) ;
    mux21_ni ix113 (.Y (sub_value[13]), .A0 (Adder2_value_13), .A1 (
             Adder1_value_13), .S0 (nx456)) ;
    mux21_ni ix121 (.Y (sub_value[14]), .A0 (Adder2_value_14), .A1 (
             Adder1_value_14), .S0 (nx456)) ;
    mux21_ni ix129 (.Y (sub_value[15]), .A0 (Adder2_value_15), .A1 (
             Adder1_value_15), .S0 (nx456)) ;
    nor02ii ix1 (.Y (sub_value[16]), .A0 (nx456), .A1 (Adder2_value_16)) ;
    mux21_ni ix137 (.Y (sub_value[17]), .A0 (Adder2_value_17), .A1 (
             Adder1_value_17), .S0 (nx456)) ;
    inv02 ix451 (.Y (nx452), .A (Adder1_value_16)) ;
    inv02 ix453 (.Y (nx454), .A (Adder1_value_16)) ;
    inv02 ix455 (.Y (nx456), .A (Adder1_value_16)) ;
endmodule


module nbit_adder_18 ( a, b, cin, add_out ) ;

    input [17:0]a ;
    input [17:0]b ;
    input cin ;
    output [17:0]add_out ;

    wire temp_16, temp_15, temp_14, temp_13, temp_12, temp_11, temp_10, temp_9, 
         temp_8, temp_7, temp_6, temp_5, temp_4, temp_3, temp_2, temp_1, temp_0;
    wire [0:0] \$dummy ;




    bit_adder f0 (.a (a[0]), .b (b[0]), .cin (cin), .s (add_out[0]), .cout (
              temp_0)) ;
    bit_adder loop1_1_fx (.a (a[1]), .b (b[1]), .cin (temp_0), .s (add_out[1]), 
              .cout (temp_1)) ;
    bit_adder loop1_2_fx (.a (a[2]), .b (b[2]), .cin (temp_1), .s (add_out[2]), 
              .cout (temp_2)) ;
    bit_adder loop1_3_fx (.a (a[3]), .b (b[3]), .cin (temp_2), .s (add_out[3]), 
              .cout (temp_3)) ;
    bit_adder loop1_4_fx (.a (a[4]), .b (b[4]), .cin (temp_3), .s (add_out[4]), 
              .cout (temp_4)) ;
    bit_adder loop1_5_fx (.a (a[5]), .b (b[5]), .cin (temp_4), .s (add_out[5]), 
              .cout (temp_5)) ;
    bit_adder loop1_6_fx (.a (a[6]), .b (b[6]), .cin (temp_5), .s (add_out[6]), 
              .cout (temp_6)) ;
    bit_adder loop1_7_fx (.a (a[7]), .b (b[7]), .cin (temp_6), .s (add_out[7]), 
              .cout (temp_7)) ;
    bit_adder loop1_8_fx (.a (a[8]), .b (b[8]), .cin (temp_7), .s (add_out[8]), 
              .cout (temp_8)) ;
    bit_adder loop1_9_fx (.a (a[9]), .b (b[9]), .cin (temp_8), .s (add_out[9]), 
              .cout (temp_9)) ;
    bit_adder loop1_10_fx (.a (a[10]), .b (b[10]), .cin (temp_9), .s (
              add_out[10]), .cout (temp_10)) ;
    bit_adder loop1_11_fx (.a (a[11]), .b (b[11]), .cin (temp_10), .s (
              add_out[11]), .cout (temp_11)) ;
    bit_adder loop1_12_fx (.a (a[12]), .b (b[12]), .cin (temp_11), .s (
              add_out[12]), .cout (temp_12)) ;
    bit_adder loop1_13_fx (.a (a[13]), .b (b[13]), .cin (temp_12), .s (
              add_out[13]), .cout (temp_13)) ;
    bit_adder loop1_14_fx (.a (a[14]), .b (b[14]), .cin (temp_13), .s (
              add_out[14]), .cout (temp_14)) ;
    bit_adder loop1_15_fx (.a (a[15]), .b (b[15]), .cin (temp_14), .s (
              add_out[15]), .cout (temp_15)) ;
    bit_adder loop1_16_fx (.a (a[16]), .b (b[16]), .cin (temp_15), .s (
              add_out[16]), .cout (temp_16)) ;
    bit_adder loop1_17_fx (.a (a[17]), .b (b[17]), .cin (temp_16), .s (
              add_out[17]), .cout (\$dummy [0])) ;
endmodule


module bit_adder ( a, b, cin, s, cout ) ;

    input a ;
    input b ;
    input cin ;
    output s ;
    output cout ;

    wire nx0, nx109;



    ao22 ix7 (.Y (cout), .A0 (b), .A1 (a), .B0 (cin), .B1 (nx0)) ;
    xnor2 ix9 (.Y (s), .A0 (nx109), .A1 (cin)) ;
    xnor2 ix110 (.Y (nx109), .A0 (a), .A1 (b)) ;
    inv01 ix1 (.Y (nx0), .A (nx109)) ;
endmodule


module selectData ( inc_dec, s, address, func ) ;

    input inc_dec ;
    input [1:0]s ;
    input [7:0]address ;
    output func ;

    wire nx12, nx38, nx52, nx72, nx181, nx183, nx186, nx188, nx191, nx193, nx195, 
         nx197;



    mux21_ni ix77 (.Y (func), .A0 (nx38), .A1 (nx72), .S0 (s[0])) ;
    nand03 ix39 (.Y (nx38), .A0 (nx181), .A1 (s[1]), .A2 (nx186)) ;
    nand02 ix182 (.Y (nx181), .A0 (nx183), .A1 (nx12)) ;
    inv01 ix184 (.Y (nx183), .A (inc_dec)) ;
    nor04 ix13 (.Y (nx12), .A0 (address[7]), .A1 (address[6]), .A2 (address[5])
          , .A3 (address[4])) ;
    mux21_ni ix187 (.Y (nx186), .A0 (nx183), .A1 (nx12), .S0 (nx188)) ;
    nand04 ix189 (.Y (nx188), .A0 (address[7]), .A1 (address[6]), .A2 (
           address[5]), .A3 (address[4])) ;
    nand03 ix73 (.Y (nx72), .A0 (nx191), .A1 (nx195), .A2 (nx197)) ;
    mux21_ni ix192 (.Y (nx191), .A0 (nx193), .A1 (address[2]), .S0 (address[1])
             ) ;
    inv01 ix194 (.Y (nx193), .A (address[0])) ;
    inv01 ix196 (.Y (nx195), .A (s[1])) ;
    aoi221 ix198 (.Y (nx197), .A0 (address[2]), .A1 (inc_dec), .B0 (address[3])
           , .B1 (nx193), .C0 (nx52)) ;
    nor02_2x ix53 (.Y (nx52), .A0 (address[3]), .A1 (inc_dec)) ;
endmodule


module nbit_mux3x1_8 ( input1, input2, input3, s, \output  ) ;

    input [7:0]input1 ;
    input [7:0]input2 ;
    input [7:0]input3 ;
    input [1:0]s ;
    output [7:0]\output  ;

    wire nx4, nx12, nx100, nx105, nx108, nx111, nx114, nx117, nx120, nx123, 
         nx130, nx132, nx134, nx140, nx142;



    inv01 ix19 (.Y (\output [0]), .A (nx100)) ;
    aoi222 ix101 (.Y (nx100), .A0 (input3[0]), .A1 (nx140), .B0 (input1[0]), .B1 (
           nx134), .C0 (input2[0]), .C1 (nx130)) ;
    nor02_2x ix13 (.Y (nx12), .A0 (nx140), .A1 (s[0])) ;
    nor02ii ix5 (.Y (nx4), .A0 (nx140), .A1 (s[0])) ;
    inv01 ix29 (.Y (\output [1]), .A (nx105)) ;
    aoi222 ix106 (.Y (nx105), .A0 (input3[1]), .A1 (nx140), .B0 (input1[1]), .B1 (
           nx134), .C0 (input2[1]), .C1 (nx130)) ;
    inv01 ix39 (.Y (\output [2]), .A (nx108)) ;
    aoi222 ix109 (.Y (nx108), .A0 (input3[2]), .A1 (nx140), .B0 (input1[2]), .B1 (
           nx134), .C0 (input2[2]), .C1 (nx130)) ;
    inv01 ix49 (.Y (\output [3]), .A (nx111)) ;
    aoi222 ix112 (.Y (nx111), .A0 (input3[3]), .A1 (nx140), .B0 (input1[3]), .B1 (
           nx134), .C0 (input2[3]), .C1 (nx130)) ;
    inv01 ix59 (.Y (\output [4]), .A (nx114)) ;
    aoi222 ix115 (.Y (nx114), .A0 (input3[4]), .A1 (nx140), .B0 (input1[4]), .B1 (
           nx134), .C0 (input2[4]), .C1 (nx130)) ;
    inv01 ix69 (.Y (\output [5]), .A (nx117)) ;
    aoi222 ix118 (.Y (nx117), .A0 (input3[5]), .A1 (nx142), .B0 (input1[5]), .B1 (
           nx134), .C0 (input2[5]), .C1 (nx130)) ;
    inv01 ix79 (.Y (\output [6]), .A (nx120)) ;
    aoi222 ix121 (.Y (nx120), .A0 (input3[6]), .A1 (nx142), .B0 (input1[6]), .B1 (
           nx12), .C0 (input2[6]), .C1 (nx130)) ;
    inv01 ix89 (.Y (\output [7]), .A (nx123)) ;
    aoi222 ix124 (.Y (nx123), .A0 (nx142), .A1 (input3[7]), .B0 (input1[7]), .B1 (
           nx12), .C0 (input2[7]), .C1 (nx132)) ;
    buf02 ix129 (.Y (nx130), .A (nx4)) ;
    buf02 ix131 (.Y (nx132), .A (nx4)) ;
    nor02_2x ix133 (.Y (nx134), .A0 (nx142), .A1 (s[0])) ;
    buf02 ix139 (.Y (nx140), .A (s[1])) ;
    buf02 ix141 (.Y (nx142), .A (s[1])) ;
endmodule


module nbit_Register_1 ( Clk, rst, enable, d, rst_value, q ) ;

    input Clk ;
    input rst ;
    input enable ;
    input [0:0]d ;
    input [0:0]rst_value ;
    output [0:0]q ;

    wire nx8, nx77, nx90;
    wire [0:0] \$dummy ;




    dff reg_q_0 (.Q (q[0]), .QB (\$dummy [0]), .D (nx77), .CLK (Clk)) ;
    mux21_ni ix78 (.Y (nx77), .A0 (nx8), .A1 (q[0]), .S0 (nx90)) ;
    mux21_ni ix9 (.Y (nx8), .A0 (d[0]), .A1 (rst_value[0]), .S0 (rst)) ;
    nor02_2x ix91 (.Y (nx90), .A0 (rst), .A1 (enable)) ;
endmodule


module nbit_Register_12 ( Clk, rst, enable, d, rst_value, q ) ;

    input Clk ;
    input rst ;
    input enable ;
    input [11:0]d ;
    input [11:0]rst_value ;
    output [11:0]q ;

    wire nx8, nx22, nx36, nx50, nx64, nx78, nx92, nx106, nx120, nx134, nx148, 
         nx162, nx286, nx296, nx306, nx316, nx326, nx336, nx346, nx356, nx366, 
         nx376, nx386, nx396, nx409, nx461, nx467, nx469;
    wire [11:0] \$dummy ;




    dff reg_q_0 (.Q (q[0]), .QB (\$dummy [0]), .D (nx286), .CLK (Clk)) ;
    mux21_ni ix287 (.Y (nx286), .A0 (nx8), .A1 (q[0]), .S0 (nx461)) ;
    mux21_ni ix9 (.Y (nx8), .A0 (d[0]), .A1 (rst_value[0]), .S0 (nx467)) ;
    nor02_2x ix410 (.Y (nx409), .A0 (nx467), .A1 (enable)) ;
    dff reg_q_1 (.Q (q[1]), .QB (\$dummy [1]), .D (nx296), .CLK (Clk)) ;
    mux21_ni ix297 (.Y (nx296), .A0 (nx22), .A1 (q[1]), .S0 (nx461)) ;
    mux21_ni ix23 (.Y (nx22), .A0 (d[1]), .A1 (rst_value[1]), .S0 (nx467)) ;
    dff reg_q_2 (.Q (q[2]), .QB (\$dummy [2]), .D (nx306), .CLK (Clk)) ;
    mux21_ni ix307 (.Y (nx306), .A0 (nx36), .A1 (q[2]), .S0 (nx461)) ;
    mux21_ni ix37 (.Y (nx36), .A0 (d[2]), .A1 (rst_value[2]), .S0 (nx467)) ;
    dff reg_q_3 (.Q (q[3]), .QB (\$dummy [3]), .D (nx316), .CLK (Clk)) ;
    mux21_ni ix317 (.Y (nx316), .A0 (nx50), .A1 (q[3]), .S0 (nx461)) ;
    mux21_ni ix51 (.Y (nx50), .A0 (d[3]), .A1 (rst_value[3]), .S0 (nx467)) ;
    dff reg_q_4 (.Q (q[4]), .QB (\$dummy [4]), .D (nx326), .CLK (Clk)) ;
    mux21_ni ix327 (.Y (nx326), .A0 (nx64), .A1 (q[4]), .S0 (nx461)) ;
    mux21_ni ix65 (.Y (nx64), .A0 (d[4]), .A1 (rst_value[4]), .S0 (nx467)) ;
    dff reg_q_5 (.Q (q[5]), .QB (\$dummy [5]), .D (nx336), .CLK (Clk)) ;
    mux21_ni ix337 (.Y (nx336), .A0 (nx78), .A1 (q[5]), .S0 (nx461)) ;
    mux21_ni ix79 (.Y (nx78), .A0 (d[5]), .A1 (rst_value[5]), .S0 (nx467)) ;
    dff reg_q_6 (.Q (q[6]), .QB (\$dummy [6]), .D (nx346), .CLK (Clk)) ;
    mux21_ni ix347 (.Y (nx346), .A0 (nx92), .A1 (q[6]), .S0 (nx409)) ;
    mux21_ni ix93 (.Y (nx92), .A0 (d[6]), .A1 (rst_value[6]), .S0 (nx469)) ;
    dff reg_q_7 (.Q (q[7]), .QB (\$dummy [7]), .D (nx356), .CLK (Clk)) ;
    mux21_ni ix357 (.Y (nx356), .A0 (nx106), .A1 (q[7]), .S0 (nx409)) ;
    mux21_ni ix107 (.Y (nx106), .A0 (d[7]), .A1 (rst_value[7]), .S0 (nx469)) ;
    dff reg_q_8 (.Q (q[8]), .QB (\$dummy [8]), .D (nx366), .CLK (Clk)) ;
    mux21_ni ix367 (.Y (nx366), .A0 (nx120), .A1 (q[8]), .S0 (nx409)) ;
    mux21_ni ix121 (.Y (nx120), .A0 (d[8]), .A1 (rst_value[8]), .S0 (nx469)) ;
    dff reg_q_9 (.Q (q[9]), .QB (\$dummy [9]), .D (nx376), .CLK (Clk)) ;
    mux21_ni ix377 (.Y (nx376), .A0 (nx134), .A1 (q[9]), .S0 (nx409)) ;
    mux21_ni ix135 (.Y (nx134), .A0 (d[9]), .A1 (rst_value[9]), .S0 (nx469)) ;
    dff reg_q_10 (.Q (q[10]), .QB (\$dummy [10]), .D (nx386), .CLK (Clk)) ;
    mux21_ni ix387 (.Y (nx386), .A0 (nx148), .A1 (q[10]), .S0 (nx409)) ;
    mux21_ni ix149 (.Y (nx148), .A0 (d[10]), .A1 (rst_value[10]), .S0 (nx469)) ;
    dff reg_q_11 (.Q (q[11]), .QB (\$dummy [11]), .D (nx396), .CLK (Clk)) ;
    mux21_ni ix397 (.Y (nx396), .A0 (nx162), .A1 (q[11]), .S0 (nx409)) ;
    mux21_ni ix163 (.Y (nx162), .A0 (d[11]), .A1 (rst_value[11]), .S0 (nx469)) ;
    nor02_2x ix460 (.Y (nx461), .A0 (nx469), .A1 (enable)) ;
    buf02 ix466 (.Y (nx467), .A (rst)) ;
    buf02 ix468 (.Y (nx469), .A (rst)) ;
endmodule


module nbit_Register_8 ( Clk, rst, enable, d, rst_value, q ) ;

    input Clk ;
    input rst ;
    input enable ;
    input [7:0]d ;
    input [7:0]rst_value ;
    output [7:0]q ;

    wire nx8, nx22, nx36, nx50, nx64, nx78, nx92, nx106, nx210, nx220, nx230, 
         nx240, nx250, nx260, nx270, nx280, nx293, nx329, nx335, nx337;
    wire [7:0] \$dummy ;




    dff reg_q_0 (.Q (q[0]), .QB (\$dummy [0]), .D (nx210), .CLK (Clk)) ;
    mux21_ni ix211 (.Y (nx210), .A0 (nx8), .A1 (q[0]), .S0 (nx329)) ;
    mux21_ni ix9 (.Y (nx8), .A0 (d[0]), .A1 (rst_value[0]), .S0 (nx335)) ;
    nor02_2x ix294 (.Y (nx293), .A0 (nx335), .A1 (enable)) ;
    dff reg_q_1 (.Q (q[1]), .QB (\$dummy [1]), .D (nx220), .CLK (Clk)) ;
    mux21_ni ix221 (.Y (nx220), .A0 (nx22), .A1 (q[1]), .S0 (nx329)) ;
    mux21_ni ix23 (.Y (nx22), .A0 (d[1]), .A1 (rst_value[1]), .S0 (nx335)) ;
    dff reg_q_2 (.Q (q[2]), .QB (\$dummy [2]), .D (nx230), .CLK (Clk)) ;
    mux21_ni ix231 (.Y (nx230), .A0 (nx36), .A1 (q[2]), .S0 (nx329)) ;
    mux21_ni ix37 (.Y (nx36), .A0 (d[2]), .A1 (rst_value[2]), .S0 (nx335)) ;
    dff reg_q_3 (.Q (q[3]), .QB (\$dummy [3]), .D (nx240), .CLK (Clk)) ;
    mux21_ni ix241 (.Y (nx240), .A0 (nx50), .A1 (q[3]), .S0 (nx329)) ;
    mux21_ni ix51 (.Y (nx50), .A0 (d[3]), .A1 (rst_value[3]), .S0 (nx335)) ;
    dff reg_q_4 (.Q (q[4]), .QB (\$dummy [4]), .D (nx250), .CLK (Clk)) ;
    mux21_ni ix251 (.Y (nx250), .A0 (nx64), .A1 (q[4]), .S0 (nx329)) ;
    mux21_ni ix65 (.Y (nx64), .A0 (d[4]), .A1 (rst_value[4]), .S0 (nx335)) ;
    dff reg_q_5 (.Q (q[5]), .QB (\$dummy [5]), .D (nx260), .CLK (Clk)) ;
    mux21_ni ix261 (.Y (nx260), .A0 (nx78), .A1 (q[5]), .S0 (nx329)) ;
    mux21_ni ix79 (.Y (nx78), .A0 (d[5]), .A1 (rst_value[5]), .S0 (nx335)) ;
    dff reg_q_6 (.Q (q[6]), .QB (\$dummy [6]), .D (nx270), .CLK (Clk)) ;
    mux21_ni ix271 (.Y (nx270), .A0 (nx92), .A1 (q[6]), .S0 (nx293)) ;
    mux21_ni ix93 (.Y (nx92), .A0 (d[6]), .A1 (rst_value[6]), .S0 (nx337)) ;
    dff reg_q_7 (.Q (q[7]), .QB (\$dummy [7]), .D (nx280), .CLK (Clk)) ;
    mux21_ni ix281 (.Y (nx280), .A0 (nx106), .A1 (q[7]), .S0 (nx293)) ;
    mux21_ni ix107 (.Y (nx106), .A0 (d[7]), .A1 (rst_value[7]), .S0 (nx337)) ;
    nor02_2x ix328 (.Y (nx329), .A0 (nx337), .A1 (enable)) ;
    buf02 ix334 (.Y (nx335), .A (rst)) ;
    buf02 ix336 (.Y (nx337), .A (rst)) ;
endmodule


module nbit_Register_18 ( Clk, rst, enable, d, rst_value, q ) ;

    input Clk ;
    input rst ;
    input enable ;
    input [17:0]d ;
    input [17:0]rst_value ;
    output [17:0]q ;

    wire nx8, nx22, nx36, nx50, nx64, nx78, nx92, nx106, nx120, nx134, nx148, 
         nx162, nx176, nx190, nx204, nx218, nx232, nx246, nx400, nx410, nx420, 
         nx430, nx440, nx450, nx460, nx470, nx480, nx490, nx500, nx510, nx520, 
         nx530, nx540, nx550, nx560, nx570, nx583, nx659, nx661, nx667, nx669, 
         nx671, nx673;
    wire [17:0] \$dummy ;




    dff reg_q_0 (.Q (q[0]), .QB (\$dummy [0]), .D (nx400), .CLK (Clk)) ;
    mux21_ni ix401 (.Y (nx400), .A0 (nx8), .A1 (q[0]), .S0 (nx659)) ;
    mux21_ni ix9 (.Y (nx8), .A0 (d[0]), .A1 (rst_value[0]), .S0 (nx669)) ;
    nor02_2x ix584 (.Y (nx583), .A0 (nx669), .A1 (enable)) ;
    dff reg_q_1 (.Q (q[1]), .QB (\$dummy [1]), .D (nx410), .CLK (Clk)) ;
    mux21_ni ix411 (.Y (nx410), .A0 (nx22), .A1 (q[1]), .S0 (nx659)) ;
    mux21_ni ix23 (.Y (nx22), .A0 (d[1]), .A1 (rst_value[1]), .S0 (nx669)) ;
    dff reg_q_2 (.Q (q[2]), .QB (\$dummy [2]), .D (nx420), .CLK (Clk)) ;
    mux21_ni ix421 (.Y (nx420), .A0 (nx36), .A1 (q[2]), .S0 (nx659)) ;
    mux21_ni ix37 (.Y (nx36), .A0 (d[2]), .A1 (rst_value[2]), .S0 (nx669)) ;
    dff reg_q_3 (.Q (q[3]), .QB (\$dummy [3]), .D (nx430), .CLK (Clk)) ;
    mux21_ni ix431 (.Y (nx430), .A0 (nx50), .A1 (q[3]), .S0 (nx659)) ;
    mux21_ni ix51 (.Y (nx50), .A0 (d[3]), .A1 (rst_value[3]), .S0 (nx669)) ;
    dff reg_q_4 (.Q (q[4]), .QB (\$dummy [4]), .D (nx440), .CLK (Clk)) ;
    mux21_ni ix441 (.Y (nx440), .A0 (nx64), .A1 (q[4]), .S0 (nx659)) ;
    mux21_ni ix65 (.Y (nx64), .A0 (d[4]), .A1 (rst_value[4]), .S0 (nx669)) ;
    dff reg_q_5 (.Q (q[5]), .QB (\$dummy [5]), .D (nx450), .CLK (Clk)) ;
    mux21_ni ix451 (.Y (nx450), .A0 (nx78), .A1 (q[5]), .S0 (nx659)) ;
    mux21_ni ix79 (.Y (nx78), .A0 (d[5]), .A1 (rst_value[5]), .S0 (nx669)) ;
    dff reg_q_6 (.Q (q[6]), .QB (\$dummy [6]), .D (nx460), .CLK (Clk)) ;
    mux21_ni ix461 (.Y (nx460), .A0 (nx92), .A1 (q[6]), .S0 (nx661)) ;
    mux21_ni ix93 (.Y (nx92), .A0 (d[6]), .A1 (rst_value[6]), .S0 (nx671)) ;
    dff reg_q_7 (.Q (q[7]), .QB (\$dummy [7]), .D (nx470), .CLK (Clk)) ;
    mux21_ni ix471 (.Y (nx470), .A0 (nx106), .A1 (q[7]), .S0 (nx661)) ;
    mux21_ni ix107 (.Y (nx106), .A0 (d[7]), .A1 (rst_value[7]), .S0 (nx671)) ;
    dff reg_q_8 (.Q (q[8]), .QB (\$dummy [8]), .D (nx480), .CLK (Clk)) ;
    mux21_ni ix481 (.Y (nx480), .A0 (nx120), .A1 (q[8]), .S0 (nx661)) ;
    mux21_ni ix121 (.Y (nx120), .A0 (d[8]), .A1 (rst_value[8]), .S0 (nx671)) ;
    dff reg_q_9 (.Q (q[9]), .QB (\$dummy [9]), .D (nx490), .CLK (Clk)) ;
    mux21_ni ix491 (.Y (nx490), .A0 (nx134), .A1 (q[9]), .S0 (nx661)) ;
    mux21_ni ix135 (.Y (nx134), .A0 (d[9]), .A1 (rst_value[9]), .S0 (nx671)) ;
    dff reg_q_10 (.Q (q[10]), .QB (\$dummy [10]), .D (nx500), .CLK (Clk)) ;
    mux21_ni ix501 (.Y (nx500), .A0 (nx148), .A1 (q[10]), .S0 (nx661)) ;
    mux21_ni ix149 (.Y (nx148), .A0 (d[10]), .A1 (rst_value[10]), .S0 (nx671)) ;
    dff reg_q_11 (.Q (q[11]), .QB (\$dummy [11]), .D (nx510), .CLK (Clk)) ;
    mux21_ni ix511 (.Y (nx510), .A0 (nx162), .A1 (q[11]), .S0 (nx661)) ;
    mux21_ni ix163 (.Y (nx162), .A0 (d[11]), .A1 (rst_value[11]), .S0 (nx671)) ;
    dff reg_q_12 (.Q (q[12]), .QB (\$dummy [12]), .D (nx520), .CLK (Clk)) ;
    mux21_ni ix521 (.Y (nx520), .A0 (nx176), .A1 (q[12]), .S0 (nx583)) ;
    mux21_ni ix177 (.Y (nx176), .A0 (d[12]), .A1 (rst_value[12]), .S0 (nx671)) ;
    dff reg_q_13 (.Q (q[13]), .QB (\$dummy [13]), .D (nx530), .CLK (Clk)) ;
    mux21_ni ix531 (.Y (nx530), .A0 (nx190), .A1 (q[13]), .S0 (nx583)) ;
    mux21_ni ix191 (.Y (nx190), .A0 (d[13]), .A1 (rst_value[13]), .S0 (nx673)) ;
    dff reg_q_14 (.Q (q[14]), .QB (\$dummy [14]), .D (nx540), .CLK (Clk)) ;
    mux21_ni ix541 (.Y (nx540), .A0 (nx204), .A1 (q[14]), .S0 (nx583)) ;
    mux21_ni ix205 (.Y (nx204), .A0 (d[14]), .A1 (rst_value[14]), .S0 (nx673)) ;
    dff reg_q_15 (.Q (q[15]), .QB (\$dummy [15]), .D (nx550), .CLK (Clk)) ;
    mux21_ni ix551 (.Y (nx550), .A0 (nx218), .A1 (q[15]), .S0 (nx583)) ;
    mux21_ni ix219 (.Y (nx218), .A0 (d[15]), .A1 (rst_value[15]), .S0 (nx673)) ;
    dff reg_q_16 (.Q (q[16]), .QB (\$dummy [16]), .D (nx560), .CLK (Clk)) ;
    mux21_ni ix561 (.Y (nx560), .A0 (nx232), .A1 (q[16]), .S0 (nx583)) ;
    mux21_ni ix233 (.Y (nx232), .A0 (d[16]), .A1 (rst_value[16]), .S0 (nx673)) ;
    dff reg_q_17 (.Q (q[17]), .QB (\$dummy [17]), .D (nx570), .CLK (Clk)) ;
    mux21_ni ix571 (.Y (nx570), .A0 (nx246), .A1 (q[17]), .S0 (nx583)) ;
    mux21_ni ix247 (.Y (nx246), .A0 (d[17]), .A1 (rst_value[17]), .S0 (nx673)) ;
    nor02_2x ix658 (.Y (nx659), .A0 (nx673), .A1 (enable)) ;
    nor02_2x ix660 (.Y (nx661), .A0 (nx673), .A1 (enable)) ;
    inv01 ix666 (.Y (nx667), .A (rst)) ;
    inv02 ix668 (.Y (nx669), .A (nx667)) ;
    inv02 ix670 (.Y (nx671), .A (nx667)) ;
    inv02 ix672 (.Y (nx673), .A (nx667)) ;
endmodule


module CacheMemory ( clk, rst, write_en, address, datain, dataout ) ;

    input clk ;
    input rst ;
    input write_en ;
    input [7:0]address ;
    input [7:0]datain ;
    output [7:0]dataout ;

    wire nx10, ram_191__0, nx24, nx32, ram_190__0, nx46, nx54, ram_189__0, nx70, 
         nx78, ram_188__0, nx90, nx98, ram_187__0, nx116, nx124, ram_186__0, 
         nx134, nx142, ram_185__0, nx154, nx162, ram_184__0, nx172, nx180, nx194, 
         ram_183__0, nx200, nx208, ram_182__0, nx218, nx226, ram_181__0, nx238, 
         nx246, ram_180__0, nx256, nx264, ram_179__0, nx280, nx288, ram_178__0, 
         nx298, nx306, ram_177__0, nx318, nx326, ram_176__0, nx344, nx358, nx370, 
         ram_175__0, nx378, ram_174__0, nx394, ram_173__0, nx412, ram_172__0, 
         nx428, ram_171__0, nx448, ram_170__0, nx464, ram_169__0, nx482, 
         ram_168__0, nx498, nx512, ram_167__0, nx520, ram_166__0, nx536, 
         ram_165__0, nx554, ram_164__0, nx570, ram_163__0, nx590, ram_162__0, 
         nx606, ram_161__0, nx624, ram_160__0, nx640, nx654, nx668, ram_159__0, 
         nx676, ram_158__0, nx692, ram_157__0, nx710, ram_156__0, nx726, 
         ram_155__0, nx746, ram_154__0, nx762, ram_153__0, nx780, ram_152__0, 
         nx796, nx810, ram_151__0, nx818, ram_150__0, nx834, ram_149__0, nx852, 
         ram_148__0, nx868, ram_147__0, nx888, ram_146__0, nx904, ram_145__0, 
         nx922, ram_144__0, nx938, nx952, nx962, ram_143__0, nx970, ram_142__0, 
         nx986, ram_141__0, nx1004, ram_140__0, nx1020, ram_139__0, nx1040, 
         ram_138__0, nx1056, ram_137__0, nx1074, ram_136__0, nx1090, nx1104, 
         ram_135__0, nx1112, ram_134__0, nx1128, ram_133__0, nx1146, ram_132__0, 
         nx1162, ram_131__0, nx1182, ram_130__0, nx1198, ram_129__0, nx1216, 
         ram_128__0, nx1232, nx1246, nx1256, nx1262, ram_127__0, nx1270, 
         ram_126__0, nx1286, ram_125__0, nx1304, ram_124__0, nx1320, ram_123__0, 
         nx1340, ram_122__0, nx1356, ram_121__0, nx1374, ram_120__0, nx1390, 
         nx1404, ram_119__0, nx1412, ram_118__0, nx1428, ram_117__0, nx1446, 
         ram_116__0, nx1462, ram_115__0, nx1482, ram_114__0, nx1498, ram_113__0, 
         nx1516, ram_112__0, nx1532, nx1546, nx1554, ram_111__0, nx1562, 
         ram_110__0, nx1578, ram_109__0, nx1596, ram_108__0, nx1612, ram_107__0, 
         nx1632, ram_106__0, nx1648, ram_105__0, nx1666, ram_104__0, nx1682, 
         nx1696, ram_103__0, nx1704, ram_102__0, nx1720, ram_101__0, nx1738, 
         ram_100__0, nx1754, ram_99__0, nx1774, ram_98__0, nx1790, ram_97__0, 
         nx1808, ram_96__0, nx1824, nx1838, ram_15__0, ram_14__0, ram_13__0, 
         ram_12__0, ram_11__0, ram_10__0, ram_9__0, ram_8__0, nx1992, ram_7__0, 
         ram_6__0, ram_5__0, ram_4__0, ram_3__0, ram_2__0, ram_1__0, ram_0__0, 
         nx2134, nx2142, ram_31__0, nx2150, ram_30__0, nx2166, ram_29__0, nx2184, 
         ram_28__0, nx2200, ram_27__0, nx2220, ram_26__0, nx2236, ram_25__0, 
         nx2254, ram_24__0, nx2270, nx2284, ram_23__0, nx2292, ram_22__0, nx2308, 
         ram_21__0, nx2326, ram_20__0, nx2342, ram_19__0, nx2362, ram_18__0, 
         nx2378, ram_17__0, nx2396, ram_16__0, nx2412, nx2426, nx2436, nx2440, 
         ram_47__0, nx2448, ram_46__0, nx2464, ram_45__0, nx2482, ram_44__0, 
         nx2498, ram_43__0, nx2518, ram_42__0, nx2534, ram_41__0, nx2552, 
         ram_40__0, nx2568, nx2582, ram_39__0, nx2590, ram_38__0, nx2606, 
         ram_37__0, nx2624, ram_36__0, nx2640, ram_35__0, nx2660, ram_34__0, 
         nx2676, ram_33__0, nx2694, ram_32__0, nx2710, nx2724, nx2732, ram_63__0, 
         nx2740, ram_62__0, nx2756, ram_61__0, nx2774, ram_60__0, nx2790, 
         ram_59__0, nx2810, ram_58__0, nx2826, ram_57__0, nx2844, ram_56__0, 
         nx2860, nx2874, ram_55__0, nx2882, ram_54__0, nx2898, ram_53__0, nx2916, 
         ram_52__0, nx2932, ram_51__0, nx2952, ram_50__0, nx2968, ram_49__0, 
         nx2986, ram_48__0, nx3002, nx3016, nx3026, ram_79__0, nx3034, ram_78__0, 
         nx3050, ram_77__0, nx3068, ram_76__0, nx3084, ram_75__0, nx3104, 
         ram_74__0, nx3120, ram_73__0, nx3138, ram_72__0, nx3154, nx3168, 
         ram_71__0, nx3176, ram_70__0, nx3192, ram_69__0, nx3210, ram_68__0, 
         nx3226, ram_67__0, nx3246, ram_66__0, nx3262, ram_65__0, nx3280, 
         ram_64__0, nx3296, nx3310, nx3318, ram_95__0, nx3326, ram_94__0, nx3342, 
         ram_93__0, nx3360, ram_92__0, nx3376, ram_91__0, nx3396, ram_90__0, 
         nx3412, ram_89__0, nx3430, ram_88__0, nx3446, nx3460, ram_87__0, nx3468, 
         ram_86__0, nx3484, ram_85__0, nx3502, ram_84__0, nx3518, ram_83__0, 
         nx3538, ram_82__0, nx3554, ram_81__0, nx3572, ram_80__0, nx3588, nx3602, 
         nx3612, nx3620, ram_207__0, nx3628, ram_206__0, nx3644, ram_205__0, 
         nx3662, ram_204__0, nx3678, ram_203__0, nx3698, ram_202__0, nx3714, 
         ram_201__0, nx3732, ram_200__0, nx3748, nx3762, ram_199__0, nx3770, 
         ram_198__0, nx3786, ram_197__0, nx3804, ram_196__0, nx3820, ram_195__0, 
         nx3840, ram_194__0, nx3856, ram_193__0, nx3874, ram_192__0, nx3890, 
         nx3904, nx3912, ram_223__0, nx3920, ram_222__0, nx3936, ram_221__0, 
         nx3954, ram_220__0, nx3970, ram_219__0, nx3990, ram_218__0, nx4006, 
         ram_217__0, nx4024, ram_216__0, nx4040, nx4054, ram_215__0, nx4062, 
         ram_214__0, nx4078, ram_213__0, nx4096, ram_212__0, nx4112, ram_211__0, 
         nx4132, ram_210__0, nx4148, ram_209__0, nx4166, ram_208__0, nx4182, 
         nx4196, nx4206, ram_239__0, nx4214, ram_238__0, nx4230, ram_237__0, 
         nx4248, ram_236__0, nx4264, ram_235__0, nx4284, ram_234__0, nx4300, 
         ram_233__0, nx4318, ram_232__0, nx4334, nx4348, ram_231__0, nx4356, 
         ram_230__0, nx4372, ram_229__0, nx4390, ram_228__0, nx4406, ram_227__0, 
         nx4426, ram_226__0, nx4442, ram_225__0, nx4460, ram_224__0, nx4476, 
         nx4490, nx4498, ram_255__0, nx4506, ram_254__0, nx4522, ram_253__0, 
         nx4540, ram_252__0, nx4556, ram_251__0, nx4576, ram_250__0, nx4592, 
         ram_249__0, nx4610, ram_248__0, nx4626, nx4640, ram_247__0, nx4648, 
         ram_246__0, nx4664, ram_245__0, nx4682, ram_244__0, nx4698, ram_243__0, 
         nx4718, ram_242__0, nx4734, ram_241__0, nx4752, ram_240__0, nx4768, 
         nx4782, nx4792, ram_191__1, ram_190__1, ram_189__1, ram_188__1, 
         ram_187__1, ram_186__1, ram_185__1, ram_184__1, nx4874, ram_183__1, 
         ram_182__1, ram_181__1, ram_180__1, ram_179__1, ram_178__1, ram_177__1, 
         ram_176__1, nx4952, ram_175__1, ram_174__1, ram_173__1, ram_172__1, 
         ram_171__1, ram_170__1, ram_169__1, ram_168__1, nx5036, ram_167__1, 
         ram_166__1, ram_165__1, ram_164__1, ram_163__1, ram_162__1, ram_161__1, 
         ram_160__1, nx5114, ram_159__1, ram_158__1, ram_157__1, ram_156__1, 
         ram_155__1, ram_154__1, ram_153__1, ram_152__1, nx5200, ram_151__1, 
         ram_150__1, ram_149__1, ram_148__1, ram_147__1, ram_146__1, ram_145__1, 
         ram_144__1, nx5278, ram_143__1, ram_142__1, ram_141__1, ram_140__1, 
         ram_139__1, ram_138__1, ram_137__1, ram_136__1, nx5362, ram_135__1, 
         ram_134__1, ram_133__1, ram_132__1, ram_131__1, ram_130__1, ram_129__1, 
         ram_128__1, nx5440, nx5450, ram_127__1, ram_126__1, ram_125__1, 
         ram_124__1, ram_123__1, ram_122__1, ram_121__1, ram_120__1, nx5528, 
         ram_119__1, ram_118__1, ram_117__1, ram_116__1, ram_115__1, ram_114__1, 
         ram_113__1, ram_112__1, nx5606, ram_111__1, ram_110__1, ram_109__1, 
         ram_108__1, ram_107__1, ram_106__1, ram_105__1, ram_104__1, nx5690, 
         ram_103__1, ram_102__1, ram_101__1, ram_100__1, ram_99__1, ram_98__1, 
         ram_97__1, ram_96__1, nx5768, ram_15__1, ram_14__1, ram_13__1, 
         ram_12__1, ram_11__1, ram_10__1, ram_9__1, ram_8__1, nx5854, ram_7__1, 
         ram_6__1, ram_5__1, ram_4__1, ram_3__1, ram_2__1, ram_1__1, ram_0__1, 
         nx5932, ram_31__1, ram_30__1, ram_29__1, ram_28__1, ram_27__1, 
         ram_26__1, ram_25__1, ram_24__1, nx6016, ram_23__1, ram_22__1, 
         ram_21__1, ram_20__1, ram_19__1, ram_18__1, ram_17__1, ram_16__1, 
         nx6094, nx6104, ram_47__1, ram_46__1, ram_45__1, ram_44__1, ram_43__1, 
         ram_42__1, ram_41__1, ram_40__1, nx6184, ram_39__1, ram_38__1, 
         ram_37__1, ram_36__1, ram_35__1, ram_34__1, ram_33__1, ram_32__1, 
         nx6262, ram_63__1, ram_62__1, ram_61__1, ram_60__1, ram_59__1, 
         ram_58__1, ram_57__1, ram_56__1, nx6346, ram_55__1, ram_54__1, 
         ram_53__1, ram_52__1, ram_51__1, ram_50__1, ram_49__1, ram_48__1, 
         nx6424, ram_79__1, ram_78__1, ram_77__1, ram_76__1, ram_75__1, 
         ram_74__1, ram_73__1, ram_72__1, nx6510, ram_71__1, ram_70__1, 
         ram_69__1, ram_68__1, ram_67__1, ram_66__1, ram_65__1, ram_64__1, 
         nx6588, ram_95__1, ram_94__1, ram_93__1, ram_92__1, ram_91__1, 
         ram_90__1, ram_89__1, ram_88__1, nx6672, ram_87__1, ram_86__1, 
         ram_85__1, ram_84__1, ram_83__1, ram_82__1, ram_81__1, ram_80__1, 
         nx6750, nx6760, ram_207__1, ram_206__1, ram_205__1, ram_204__1, 
         ram_203__1, ram_202__1, ram_201__1, ram_200__1, nx6838, ram_199__1, 
         ram_198__1, ram_197__1, ram_196__1, ram_195__1, ram_194__1, ram_193__1, 
         ram_192__1, nx6916, ram_223__1, ram_222__1, ram_221__1, ram_220__1, 
         ram_219__1, ram_218__1, ram_217__1, ram_216__1, nx7000, ram_215__1, 
         ram_214__1, ram_213__1, ram_212__1, ram_211__1, ram_210__1, ram_209__1, 
         ram_208__1, nx7078, ram_239__1, ram_238__1, ram_237__1, ram_236__1, 
         ram_235__1, ram_234__1, ram_233__1, ram_232__1, nx7164, ram_231__1, 
         ram_230__1, ram_229__1, ram_228__1, ram_227__1, ram_226__1, ram_225__1, 
         ram_224__1, nx7242, ram_255__1, ram_254__1, ram_253__1, ram_252__1, 
         ram_251__1, ram_250__1, ram_249__1, ram_248__1, nx7326, ram_247__1, 
         ram_246__1, ram_245__1, ram_244__1, ram_243__1, ram_242__1, ram_241__1, 
         ram_240__1, nx7404, nx7414, ram_191__2, ram_190__2, ram_189__2, 
         ram_188__2, ram_187__2, ram_186__2, ram_185__2, ram_184__2, nx7496, 
         ram_183__2, ram_182__2, ram_181__2, ram_180__2, ram_179__2, ram_178__2, 
         ram_177__2, ram_176__2, nx7574, ram_175__2, ram_174__2, ram_173__2, 
         ram_172__2, ram_171__2, ram_170__2, ram_169__2, ram_168__2, nx7658, 
         ram_167__2, ram_166__2, ram_165__2, ram_164__2, ram_163__2, ram_162__2, 
         ram_161__2, ram_160__2, nx7736, ram_159__2, ram_158__2, ram_157__2, 
         ram_156__2, ram_155__2, ram_154__2, ram_153__2, ram_152__2, nx7822, 
         ram_151__2, ram_150__2, ram_149__2, ram_148__2, ram_147__2, ram_146__2, 
         ram_145__2, ram_144__2, nx7900, ram_143__2, ram_142__2, ram_141__2, 
         ram_140__2, ram_139__2, ram_138__2, ram_137__2, ram_136__2, nx7984, 
         ram_135__2, ram_134__2, ram_133__2, ram_132__2, ram_131__2, ram_130__2, 
         ram_129__2, ram_128__2, nx8062, nx8072, ram_127__2, ram_126__2, 
         ram_125__2, ram_124__2, ram_123__2, ram_122__2, ram_121__2, ram_120__2, 
         nx8150, ram_119__2, ram_118__2, ram_117__2, ram_116__2, ram_115__2, 
         ram_114__2, ram_113__2, ram_112__2, nx8228, ram_111__2, ram_110__2, 
         ram_109__2, ram_108__2, ram_107__2, ram_106__2, ram_105__2, ram_104__2, 
         nx8312, ram_103__2, ram_102__2, ram_101__2, ram_100__2, ram_99__2, 
         ram_98__2, ram_97__2, ram_96__2, nx8390, ram_15__2, ram_14__2, 
         ram_13__2, ram_12__2, ram_11__2, ram_10__2, ram_9__2, ram_8__2, nx8476, 
         ram_7__2, ram_6__2, ram_5__2, ram_4__2, ram_3__2, ram_2__2, ram_1__2, 
         ram_0__2, nx8554, ram_31__2, ram_30__2, ram_29__2, ram_28__2, ram_27__2, 
         ram_26__2, ram_25__2, ram_24__2, nx8638, ram_23__2, ram_22__2, 
         ram_21__2, ram_20__2, ram_19__2, ram_18__2, ram_17__2, ram_16__2, 
         nx8716, nx8726, ram_47__2, ram_46__2, ram_45__2, ram_44__2, ram_43__2, 
         ram_42__2, ram_41__2, ram_40__2, nx8806, ram_39__2, ram_38__2, 
         ram_37__2, ram_36__2, ram_35__2, ram_34__2, ram_33__2, ram_32__2, 
         nx8884, ram_63__2, ram_62__2, ram_61__2, ram_60__2, ram_59__2, 
         ram_58__2, ram_57__2, ram_56__2, nx8968, ram_55__2, ram_54__2, 
         ram_53__2, ram_52__2, ram_51__2, ram_50__2, ram_49__2, ram_48__2, 
         nx9046, ram_79__2, ram_78__2, ram_77__2, ram_76__2, ram_75__2, 
         ram_74__2, ram_73__2, ram_72__2, nx9132, ram_71__2, ram_70__2, 
         ram_69__2, ram_68__2, ram_67__2, ram_66__2, ram_65__2, ram_64__2, 
         nx9210, ram_95__2, ram_94__2, ram_93__2, ram_92__2, ram_91__2, 
         ram_90__2, ram_89__2, ram_88__2, nx9294, ram_87__2, ram_86__2, 
         ram_85__2, ram_84__2, ram_83__2, ram_82__2, ram_81__2, ram_80__2, 
         nx9372, nx9382, ram_207__2, ram_206__2, ram_205__2, ram_204__2, 
         ram_203__2, ram_202__2, ram_201__2, ram_200__2, nx9460, ram_199__2, 
         ram_198__2, ram_197__2, ram_196__2, ram_195__2, ram_194__2, ram_193__2, 
         ram_192__2, nx9538, ram_223__2, ram_222__2, ram_221__2, ram_220__2, 
         ram_219__2, ram_218__2, ram_217__2, ram_216__2, nx9622, ram_215__2, 
         ram_214__2, ram_213__2, ram_212__2, ram_211__2, ram_210__2, ram_209__2, 
         ram_208__2, nx9700, ram_239__2, ram_238__2, ram_237__2, ram_236__2, 
         ram_235__2, ram_234__2, ram_233__2, ram_232__2, nx9786, ram_231__2, 
         ram_230__2, ram_229__2, ram_228__2, ram_227__2, ram_226__2, ram_225__2, 
         ram_224__2, nx9864, ram_255__2, ram_254__2, ram_253__2, ram_252__2, 
         ram_251__2, ram_250__2, ram_249__2, ram_248__2, nx9948, ram_247__2, 
         ram_246__2, ram_245__2, ram_244__2, ram_243__2, ram_242__2, ram_241__2, 
         ram_240__2, nx10026, nx10036, ram_191__3, ram_190__3, ram_189__3, 
         ram_188__3, ram_187__3, ram_186__3, ram_185__3, ram_184__3, nx10118, 
         ram_183__3, ram_182__3, ram_181__3, ram_180__3, ram_179__3, ram_178__3, 
         ram_177__3, ram_176__3, nx10196, ram_175__3, ram_174__3, ram_173__3, 
         ram_172__3, ram_171__3, ram_170__3, ram_169__3, ram_168__3, nx10280, 
         ram_167__3, ram_166__3, ram_165__3, ram_164__3, ram_163__3, ram_162__3, 
         ram_161__3, ram_160__3, nx10358, ram_159__3, ram_158__3, ram_157__3, 
         ram_156__3, ram_155__3, ram_154__3, ram_153__3, ram_152__3, nx10444, 
         ram_151__3, ram_150__3, ram_149__3, ram_148__3, ram_147__3, ram_146__3, 
         ram_145__3, ram_144__3, nx10522, ram_143__3, ram_142__3, ram_141__3, 
         ram_140__3, ram_139__3, ram_138__3, ram_137__3, ram_136__3, nx10606, 
         ram_135__3, ram_134__3, ram_133__3, ram_132__3, ram_131__3, ram_130__3, 
         ram_129__3, ram_128__3, nx10684, nx10694, ram_127__3, ram_126__3, 
         ram_125__3, ram_124__3, ram_123__3, ram_122__3, ram_121__3, ram_120__3, 
         nx10772, ram_119__3, ram_118__3, ram_117__3, ram_116__3, ram_115__3, 
         ram_114__3, ram_113__3, ram_112__3, nx10850, ram_111__3, ram_110__3, 
         ram_109__3, ram_108__3, ram_107__3, ram_106__3, ram_105__3, ram_104__3, 
         nx10934, ram_103__3, ram_102__3, ram_101__3, ram_100__3, ram_99__3, 
         ram_98__3, ram_97__3, ram_96__3, nx11012, ram_15__3, ram_14__3, 
         ram_13__3, ram_12__3, ram_11__3, ram_10__3, ram_9__3, ram_8__3, nx11098, 
         ram_7__3, ram_6__3, ram_5__3, ram_4__3, ram_3__3, ram_2__3, ram_1__3, 
         ram_0__3, nx11176, ram_31__3, ram_30__3, ram_29__3, ram_28__3, 
         ram_27__3, ram_26__3, ram_25__3, ram_24__3, nx11260, ram_23__3, 
         ram_22__3, ram_21__3, ram_20__3, ram_19__3, ram_18__3, ram_17__3, 
         ram_16__3, nx11338, nx11348, ram_47__3, ram_46__3, ram_45__3, ram_44__3, 
         ram_43__3, ram_42__3, ram_41__3, ram_40__3, nx11428, ram_39__3, 
         ram_38__3, ram_37__3, ram_36__3, ram_35__3, ram_34__3, ram_33__3, 
         ram_32__3, nx11506, ram_63__3, ram_62__3, ram_61__3, ram_60__3, 
         ram_59__3, ram_58__3, ram_57__3, ram_56__3, nx11590, ram_55__3, 
         ram_54__3, ram_53__3, ram_52__3, ram_51__3, ram_50__3, ram_49__3, 
         ram_48__3, nx11668, ram_79__3, ram_78__3, ram_77__3, ram_76__3, 
         ram_75__3, ram_74__3, ram_73__3, ram_72__3, nx11754, ram_71__3, 
         ram_70__3, ram_69__3, ram_68__3, ram_67__3, ram_66__3, ram_65__3, 
         ram_64__3, nx11832, ram_95__3, ram_94__3, ram_93__3, ram_92__3, 
         ram_91__3, ram_90__3, ram_89__3, ram_88__3, nx11916, ram_87__3, 
         ram_86__3, ram_85__3, ram_84__3, ram_83__3, ram_82__3, ram_81__3, 
         ram_80__3, nx11994, nx12004, ram_207__3, ram_206__3, ram_205__3, 
         ram_204__3, ram_203__3, ram_202__3, ram_201__3, ram_200__3, nx12082, 
         ram_199__3, ram_198__3, ram_197__3, ram_196__3, ram_195__3, ram_194__3, 
         ram_193__3, ram_192__3, nx12160, ram_223__3, ram_222__3, ram_221__3, 
         ram_220__3, ram_219__3, ram_218__3, ram_217__3, ram_216__3, nx12244, 
         ram_215__3, ram_214__3, ram_213__3, ram_212__3, ram_211__3, ram_210__3, 
         ram_209__3, ram_208__3, nx12322, ram_239__3, ram_238__3, ram_237__3, 
         ram_236__3, ram_235__3, ram_234__3, ram_233__3, ram_232__3, nx12408, 
         ram_231__3, ram_230__3, ram_229__3, ram_228__3, ram_227__3, ram_226__3, 
         ram_225__3, ram_224__3, nx12486, ram_255__3, ram_254__3, ram_253__3, 
         ram_252__3, ram_251__3, ram_250__3, ram_249__3, ram_248__3, nx12570, 
         ram_247__3, ram_246__3, ram_245__3, ram_244__3, ram_243__3, ram_242__3, 
         ram_241__3, ram_240__3, nx12648, nx12658, ram_191__4, ram_190__4, 
         ram_189__4, ram_188__4, ram_187__4, ram_186__4, ram_185__4, ram_184__4, 
         nx12740, ram_183__4, ram_182__4, ram_181__4, ram_180__4, ram_179__4, 
         ram_178__4, ram_177__4, ram_176__4, nx12818, ram_175__4, ram_174__4, 
         ram_173__4, ram_172__4, ram_171__4, ram_170__4, ram_169__4, ram_168__4, 
         nx12902, ram_167__4, ram_166__4, ram_165__4, ram_164__4, ram_163__4, 
         ram_162__4, ram_161__4, ram_160__4, nx12980, ram_159__4, ram_158__4, 
         ram_157__4, ram_156__4, ram_155__4, ram_154__4, ram_153__4, ram_152__4, 
         nx13066, ram_151__4, ram_150__4, ram_149__4, ram_148__4, ram_147__4, 
         ram_146__4, ram_145__4, ram_144__4, nx13144, ram_143__4, ram_142__4, 
         ram_141__4, ram_140__4, ram_139__4, ram_138__4, ram_137__4, ram_136__4, 
         nx13228, ram_135__4, ram_134__4, ram_133__4, ram_132__4, ram_131__4, 
         ram_130__4, ram_129__4, ram_128__4, nx13306, nx13316, ram_127__4, 
         ram_126__4, ram_125__4, ram_124__4, ram_123__4, ram_122__4, ram_121__4, 
         ram_120__4, nx13394, ram_119__4, ram_118__4, ram_117__4, ram_116__4, 
         ram_115__4, ram_114__4, ram_113__4, ram_112__4, nx13472, ram_111__4, 
         ram_110__4, ram_109__4, ram_108__4, ram_107__4, ram_106__4, ram_105__4, 
         ram_104__4, nx13556, ram_103__4, ram_102__4, ram_101__4, ram_100__4, 
         ram_99__4, ram_98__4, ram_97__4, ram_96__4, nx13634, ram_15__4, 
         ram_14__4, ram_13__4, ram_12__4, ram_11__4, ram_10__4, ram_9__4, 
         ram_8__4, nx13720, ram_7__4, ram_6__4, ram_5__4, ram_4__4, ram_3__4, 
         ram_2__4, ram_1__4, ram_0__4, nx13798, ram_31__4, ram_30__4, ram_29__4, 
         ram_28__4, ram_27__4, ram_26__4, ram_25__4, ram_24__4, nx13882, 
         ram_23__4, ram_22__4, ram_21__4, ram_20__4, ram_19__4, ram_18__4, 
         ram_17__4, ram_16__4, nx13960, nx13970, ram_47__4, ram_46__4, ram_45__4, 
         ram_44__4, ram_43__4, ram_42__4, ram_41__4, ram_40__4, nx14050, 
         ram_39__4, ram_38__4, ram_37__4, ram_36__4, ram_35__4, ram_34__4, 
         ram_33__4, ram_32__4, nx14128, ram_63__4, ram_62__4, ram_61__4, 
         ram_60__4, ram_59__4, ram_58__4, ram_57__4, ram_56__4, nx14212, 
         ram_55__4, ram_54__4, ram_53__4, ram_52__4, ram_51__4, ram_50__4, 
         ram_49__4, ram_48__4, nx14290, ram_79__4, ram_78__4, ram_77__4, 
         ram_76__4, ram_75__4, ram_74__4, ram_73__4, ram_72__4, nx14376, 
         ram_71__4, ram_70__4, ram_69__4, ram_68__4, ram_67__4, ram_66__4, 
         ram_65__4, ram_64__4, nx14454, ram_95__4, ram_94__4, ram_93__4, 
         ram_92__4, ram_91__4, ram_90__4, ram_89__4, ram_88__4, nx14538, 
         ram_87__4, ram_86__4, ram_85__4, ram_84__4, ram_83__4, ram_82__4, 
         ram_81__4, ram_80__4, nx14616, nx14626, ram_207__4, ram_206__4, 
         ram_205__4, ram_204__4, ram_203__4, ram_202__4, ram_201__4, ram_200__4, 
         nx14704, ram_199__4, ram_198__4, ram_197__4, ram_196__4, ram_195__4, 
         ram_194__4, ram_193__4, ram_192__4, nx14782, ram_223__4, ram_222__4, 
         ram_221__4, ram_220__4, ram_219__4, ram_218__4, ram_217__4, ram_216__4, 
         nx14866, ram_215__4, ram_214__4, ram_213__4, ram_212__4, ram_211__4, 
         ram_210__4, ram_209__4, ram_208__4, nx14944, ram_239__4, ram_238__4, 
         ram_237__4, ram_236__4, ram_235__4, ram_234__4, ram_233__4, ram_232__4, 
         nx15030, ram_231__4, ram_230__4, ram_229__4, ram_228__4, ram_227__4, 
         ram_226__4, ram_225__4, ram_224__4, nx15108, ram_255__4, ram_254__4, 
         ram_253__4, ram_252__4, ram_251__4, ram_250__4, ram_249__4, ram_248__4, 
         nx15192, ram_247__4, ram_246__4, ram_245__4, ram_244__4, ram_243__4, 
         ram_242__4, ram_241__4, ram_240__4, nx15270, nx15280, ram_191__5, 
         ram_190__5, ram_189__5, ram_188__5, ram_187__5, ram_186__5, ram_185__5, 
         ram_184__5, nx15362, ram_183__5, ram_182__5, ram_181__5, ram_180__5, 
         ram_179__5, ram_178__5, ram_177__5, ram_176__5, nx15440, ram_175__5, 
         ram_174__5, ram_173__5, ram_172__5, ram_171__5, ram_170__5, ram_169__5, 
         ram_168__5, nx15524, ram_167__5, ram_166__5, ram_165__5, ram_164__5, 
         ram_163__5, ram_162__5, ram_161__5, ram_160__5, nx15602, ram_159__5, 
         ram_158__5, ram_157__5, ram_156__5, ram_155__5, ram_154__5, ram_153__5, 
         ram_152__5, nx15688, ram_151__5, ram_150__5, ram_149__5, ram_148__5, 
         ram_147__5, ram_146__5, ram_145__5, ram_144__5, nx15766, ram_143__5, 
         ram_142__5, ram_141__5, ram_140__5, ram_139__5, ram_138__5, ram_137__5, 
         ram_136__5, nx15850, ram_135__5, ram_134__5, ram_133__5, ram_132__5, 
         ram_131__5, ram_130__5, ram_129__5, ram_128__5, nx15928, nx15938, 
         ram_127__5, ram_126__5, ram_125__5, ram_124__5, ram_123__5, ram_122__5, 
         ram_121__5, ram_120__5, nx16016, ram_119__5, ram_118__5, ram_117__5, 
         ram_116__5, ram_115__5, ram_114__5, ram_113__5, ram_112__5, nx16094, 
         ram_111__5, ram_110__5, ram_109__5, ram_108__5, ram_107__5, ram_106__5, 
         ram_105__5, ram_104__5, nx16178, ram_103__5, ram_102__5, ram_101__5, 
         ram_100__5, ram_99__5, ram_98__5, ram_97__5, ram_96__5, nx16256, 
         ram_15__5, ram_14__5, ram_13__5, ram_12__5, ram_11__5, ram_10__5, 
         ram_9__5, ram_8__5, nx16342, ram_7__5, ram_6__5, ram_5__5, ram_4__5, 
         ram_3__5, ram_2__5, ram_1__5, ram_0__5, nx16420, ram_31__5, ram_30__5, 
         ram_29__5, ram_28__5, ram_27__5, ram_26__5, ram_25__5, ram_24__5, 
         nx16504, ram_23__5, ram_22__5, ram_21__5, ram_20__5, ram_19__5, 
         ram_18__5, ram_17__5, ram_16__5, nx16582, nx16592, ram_47__5, ram_46__5, 
         ram_45__5, ram_44__5, ram_43__5, ram_42__5, ram_41__5, ram_40__5, 
         nx16672, ram_39__5, ram_38__5, ram_37__5, ram_36__5, ram_35__5, 
         ram_34__5, ram_33__5, ram_32__5, nx16750, ram_63__5, ram_62__5, 
         ram_61__5, ram_60__5, ram_59__5, ram_58__5, ram_57__5, ram_56__5, 
         nx16834, ram_55__5, ram_54__5, ram_53__5, ram_52__5, ram_51__5, 
         ram_50__5, ram_49__5, ram_48__5, nx16912, ram_79__5, ram_78__5, 
         ram_77__5, ram_76__5, ram_75__5, ram_74__5, ram_73__5, ram_72__5, 
         nx16998, ram_71__5, ram_70__5, ram_69__5, ram_68__5, ram_67__5, 
         ram_66__5, ram_65__5, ram_64__5, nx17076, ram_95__5, ram_94__5, 
         ram_93__5, ram_92__5, ram_91__5, ram_90__5, ram_89__5, ram_88__5, 
         nx17160, ram_87__5, ram_86__5, ram_85__5, ram_84__5, ram_83__5, 
         ram_82__5, ram_81__5, ram_80__5, nx17238, nx17248, ram_207__5, 
         ram_206__5, ram_205__5, ram_204__5, ram_203__5, ram_202__5, ram_201__5, 
         ram_200__5, nx17326, ram_199__5, ram_198__5, ram_197__5, ram_196__5, 
         ram_195__5, ram_194__5, ram_193__5, ram_192__5, nx17404, ram_223__5, 
         ram_222__5, ram_221__5, ram_220__5, ram_219__5, ram_218__5, ram_217__5, 
         ram_216__5, nx17488, ram_215__5, ram_214__5, ram_213__5, ram_212__5, 
         ram_211__5, ram_210__5, ram_209__5, ram_208__5, nx17566, ram_239__5, 
         ram_238__5, ram_237__5, ram_236__5, ram_235__5, ram_234__5, ram_233__5, 
         ram_232__5, nx17652, ram_231__5, ram_230__5, ram_229__5, ram_228__5, 
         ram_227__5, ram_226__5, ram_225__5, ram_224__5, nx17730, ram_255__5, 
         ram_254__5, ram_253__5, ram_252__5, ram_251__5, ram_250__5, ram_249__5, 
         ram_248__5, nx17814, ram_247__5, ram_246__5, ram_245__5, ram_244__5, 
         ram_243__5, ram_242__5, ram_241__5, ram_240__5, nx17892, nx17902, 
         ram_191__6, ram_190__6, ram_189__6, ram_188__6, ram_187__6, ram_186__6, 
         ram_185__6, ram_184__6, nx17984, ram_183__6, ram_182__6, ram_181__6, 
         ram_180__6, ram_179__6, ram_178__6, ram_177__6, ram_176__6, nx18062, 
         ram_175__6, ram_174__6, ram_173__6, ram_172__6, ram_171__6, ram_170__6, 
         ram_169__6, ram_168__6, nx18146, ram_167__6, ram_166__6, ram_165__6, 
         ram_164__6, ram_163__6, ram_162__6, ram_161__6, ram_160__6, nx18224, 
         ram_159__6, ram_158__6, ram_157__6, ram_156__6, ram_155__6, ram_154__6, 
         ram_153__6, ram_152__6, nx18310, ram_151__6, ram_150__6, ram_149__6, 
         ram_148__6, ram_147__6, ram_146__6, ram_145__6, ram_144__6, nx18388, 
         ram_143__6, ram_142__6, ram_141__6, ram_140__6, ram_139__6, ram_138__6, 
         ram_137__6, ram_136__6, nx18472, ram_135__6, ram_134__6, ram_133__6, 
         ram_132__6, ram_131__6, ram_130__6, ram_129__6, ram_128__6, nx18550, 
         nx18560, ram_127__6, ram_126__6, ram_125__6, ram_124__6, ram_123__6, 
         ram_122__6, ram_121__6, ram_120__6, nx18638, ram_119__6, ram_118__6, 
         ram_117__6, ram_116__6, ram_115__6, ram_114__6, ram_113__6, ram_112__6, 
         nx18716, ram_111__6, ram_110__6, ram_109__6, ram_108__6, ram_107__6, 
         ram_106__6, ram_105__6, ram_104__6, nx18800, ram_103__6, ram_102__6, 
         ram_101__6, ram_100__6, ram_99__6, ram_98__6, ram_97__6, ram_96__6, 
         nx18878, ram_15__6, ram_14__6, ram_13__6, ram_12__6, ram_11__6, 
         ram_10__6, ram_9__6, ram_8__6, nx18964, ram_7__6, ram_6__6, ram_5__6, 
         ram_4__6, ram_3__6, ram_2__6, ram_1__6, ram_0__6, nx19042, ram_31__6, 
         ram_30__6, ram_29__6, ram_28__6, ram_27__6, ram_26__6, ram_25__6, 
         ram_24__6, nx19126, ram_23__6, ram_22__6, ram_21__6, ram_20__6, 
         ram_19__6, ram_18__6, ram_17__6, ram_16__6, nx19204, nx19214, ram_47__6, 
         ram_46__6, ram_45__6, ram_44__6, ram_43__6, ram_42__6, ram_41__6, 
         ram_40__6, nx19294, ram_39__6, ram_38__6, ram_37__6, ram_36__6, 
         ram_35__6, ram_34__6, ram_33__6, ram_32__6, nx19372, ram_63__6, 
         ram_62__6, ram_61__6, ram_60__6, ram_59__6, ram_58__6, ram_57__6, 
         ram_56__6, nx19456, ram_55__6, ram_54__6, ram_53__6, ram_52__6, 
         ram_51__6, ram_50__6, ram_49__6, ram_48__6, nx19534, ram_79__6, 
         ram_78__6, ram_77__6, ram_76__6, ram_75__6, ram_74__6, ram_73__6, 
         ram_72__6, nx19620, ram_71__6, ram_70__6, ram_69__6, ram_68__6, 
         ram_67__6, ram_66__6, ram_65__6, ram_64__6, nx19698, ram_95__6, 
         ram_94__6, ram_93__6, ram_92__6, ram_91__6, ram_90__6, ram_89__6, 
         ram_88__6, nx19782, ram_87__6, ram_86__6, ram_85__6, ram_84__6, 
         ram_83__6, ram_82__6, ram_81__6, ram_80__6, nx19860, nx19870, 
         ram_207__6, ram_206__6, ram_205__6, ram_204__6, ram_203__6, ram_202__6, 
         ram_201__6, ram_200__6, nx19948, ram_199__6, ram_198__6, ram_197__6, 
         ram_196__6, ram_195__6, ram_194__6, ram_193__6, ram_192__6, nx20026, 
         ram_223__6, ram_222__6, ram_221__6, ram_220__6, ram_219__6, ram_218__6, 
         ram_217__6, ram_216__6, nx20110, ram_215__6, ram_214__6, ram_213__6, 
         ram_212__6, ram_211__6, ram_210__6, ram_209__6, ram_208__6, nx20188, 
         ram_239__6, ram_238__6, ram_237__6, ram_236__6, ram_235__6, ram_234__6, 
         ram_233__6, ram_232__6, nx20274, ram_231__6, ram_230__6, ram_229__6, 
         ram_228__6, ram_227__6, ram_226__6, ram_225__6, ram_224__6, nx20352, 
         ram_255__6, ram_254__6, ram_253__6, ram_252__6, ram_251__6, ram_250__6, 
         ram_249__6, ram_248__6, nx20436, ram_247__6, ram_246__6, ram_245__6, 
         ram_244__6, ram_243__6, ram_242__6, ram_241__6, ram_240__6, nx20514, 
         nx20524, ram_191__7, ram_190__7, ram_189__7, ram_188__7, ram_187__7, 
         ram_186__7, ram_185__7, ram_184__7, nx20606, ram_183__7, ram_182__7, 
         ram_181__7, ram_180__7, ram_179__7, ram_178__7, ram_177__7, ram_176__7, 
         nx20684, ram_175__7, ram_174__7, ram_173__7, ram_172__7, ram_171__7, 
         ram_170__7, ram_169__7, ram_168__7, nx20768, ram_167__7, ram_166__7, 
         ram_165__7, ram_164__7, ram_163__7, ram_162__7, ram_161__7, ram_160__7, 
         nx20846, ram_159__7, ram_158__7, ram_157__7, ram_156__7, ram_155__7, 
         ram_154__7, ram_153__7, ram_152__7, nx20932, ram_151__7, ram_150__7, 
         ram_149__7, ram_148__7, ram_147__7, ram_146__7, ram_145__7, ram_144__7, 
         nx21010, ram_143__7, ram_142__7, ram_141__7, ram_140__7, ram_139__7, 
         ram_138__7, ram_137__7, ram_136__7, nx21094, ram_135__7, ram_134__7, 
         ram_133__7, ram_132__7, ram_131__7, ram_130__7, ram_129__7, ram_128__7, 
         nx21172, nx21182, ram_127__7, ram_126__7, ram_125__7, ram_124__7, 
         ram_123__7, ram_122__7, ram_121__7, ram_120__7, nx21260, ram_119__7, 
         ram_118__7, ram_117__7, ram_116__7, ram_115__7, ram_114__7, ram_113__7, 
         ram_112__7, nx21338, ram_111__7, ram_110__7, ram_109__7, ram_108__7, 
         ram_107__7, ram_106__7, ram_105__7, ram_104__7, nx21422, ram_103__7, 
         ram_102__7, ram_101__7, ram_100__7, ram_99__7, ram_98__7, ram_97__7, 
         ram_96__7, nx21500, ram_15__7, ram_14__7, ram_13__7, ram_12__7, 
         ram_11__7, ram_10__7, ram_9__7, ram_8__7, nx21586, ram_7__7, ram_6__7, 
         ram_5__7, ram_4__7, ram_3__7, ram_2__7, ram_1__7, ram_0__7, nx21664, 
         ram_31__7, ram_30__7, ram_29__7, ram_28__7, ram_27__7, ram_26__7, 
         ram_25__7, ram_24__7, nx21748, ram_23__7, ram_22__7, ram_21__7, 
         ram_20__7, ram_19__7, ram_18__7, ram_17__7, ram_16__7, nx21826, nx21836, 
         ram_47__7, ram_46__7, ram_45__7, ram_44__7, ram_43__7, ram_42__7, 
         ram_41__7, ram_40__7, nx21916, ram_39__7, ram_38__7, ram_37__7, 
         ram_36__7, ram_35__7, ram_34__7, ram_33__7, ram_32__7, nx21994, 
         ram_63__7, ram_62__7, ram_61__7, ram_60__7, ram_59__7, ram_58__7, 
         ram_57__7, ram_56__7, nx22078, ram_55__7, ram_54__7, ram_53__7, 
         ram_52__7, ram_51__7, ram_50__7, ram_49__7, ram_48__7, nx22156, 
         ram_79__7, ram_78__7, ram_77__7, ram_76__7, ram_75__7, ram_74__7, 
         ram_73__7, ram_72__7, nx22242, ram_71__7, ram_70__7, ram_69__7, 
         ram_68__7, ram_67__7, ram_66__7, ram_65__7, ram_64__7, nx22320, 
         ram_95__7, ram_94__7, ram_93__7, ram_92__7, ram_91__7, ram_90__7, 
         ram_89__7, ram_88__7, nx22404, ram_87__7, ram_86__7, ram_85__7, 
         ram_84__7, ram_83__7, ram_82__7, ram_81__7, ram_80__7, nx22482, nx22492, 
         ram_207__7, ram_206__7, ram_205__7, ram_204__7, ram_203__7, ram_202__7, 
         ram_201__7, ram_200__7, nx22570, ram_199__7, ram_198__7, ram_197__7, 
         ram_196__7, ram_195__7, ram_194__7, ram_193__7, ram_192__7, nx22648, 
         ram_223__7, ram_222__7, ram_221__7, ram_220__7, ram_219__7, ram_218__7, 
         ram_217__7, ram_216__7, nx22732, ram_215__7, ram_214__7, ram_213__7, 
         ram_212__7, ram_211__7, ram_210__7, ram_209__7, ram_208__7, nx22810, 
         ram_239__7, ram_238__7, ram_237__7, ram_236__7, ram_235__7, ram_234__7, 
         ram_233__7, ram_232__7, nx22896, ram_231__7, ram_230__7, ram_229__7, 
         ram_228__7, ram_227__7, ram_226__7, ram_225__7, ram_224__7, nx22974, 
         ram_255__7, ram_254__7, ram_253__7, ram_252__7, ram_251__7, ram_250__7, 
         ram_249__7, ram_248__7, nx23058, ram_247__7, ram_246__7, ram_245__7, 
         ram_244__7, ram_243__7, ram_242__7, ram_241__7, ram_240__7, nx23136, 
         nx23146, nx33630, nx33640, nx33650, nx33660, nx33670, nx33680, nx33690, 
         nx33700, nx33710, nx33720, nx33730, nx33740, nx33750, nx33760, nx33770, 
         nx33780, nx33790, nx33800, nx33810, nx33820, nx33830, nx33840, nx33850, 
         nx33860, nx33870, nx33880, nx33890, nx33900, nx33910, nx33920, nx33930, 
         nx33940, nx33950, nx33960, nx33970, nx33980, nx33990, nx34000, nx34010, 
         nx34020, nx34030, nx34040, nx34050, nx34060, nx34070, nx34080, nx34090, 
         nx34100, nx34110, nx34120, nx34130, nx34140, nx34150, nx34160, nx34170, 
         nx34180, nx34190, nx34200, nx34210, nx34220, nx34230, nx34240, nx34250, 
         nx34260, nx34270, nx34280, nx34290, nx34300, nx34310, nx34320, nx34330, 
         nx34340, nx34350, nx34360, nx34370, nx34380, nx34390, nx34400, nx34410, 
         nx34420, nx34430, nx34440, nx34450, nx34460, nx34470, nx34480, nx34490, 
         nx34500, nx34510, nx34520, nx34530, nx34540, nx34550, nx34560, nx34570, 
         nx34580, nx34590, nx34600, nx34610, nx34620, nx34630, nx34640, nx34650, 
         nx34660, nx34670, nx34680, nx34690, nx34700, nx34710, nx34720, nx34730, 
         nx34740, nx34750, nx34760, nx34770, nx34780, nx34790, nx34800, nx34810, 
         nx34820, nx34830, nx34840, nx34850, nx34860, nx34870, nx34880, nx34890, 
         nx34900, nx34910, nx34920, nx34930, nx34940, nx34950, nx34960, nx34970, 
         nx34980, nx34990, nx35000, nx35010, nx35020, nx35030, nx35040, nx35050, 
         nx35060, nx35070, nx35080, nx35090, nx35100, nx35110, nx35120, nx35130, 
         nx35140, nx35150, nx35160, nx35170, nx35180, nx35190, nx35200, nx35210, 
         nx35220, nx35230, nx35240, nx35250, nx35260, nx35270, nx35280, nx35290, 
         nx35300, nx35310, nx35320, nx35330, nx35340, nx35350, nx35360, nx35370, 
         nx35380, nx35390, nx35400, nx35410, nx35420, nx35430, nx35440, nx35450, 
         nx35460, nx35470, nx35480, nx35490, nx35500, nx35510, nx35520, nx35530, 
         nx35540, nx35550, nx35560, nx35570, nx35580, nx35590, nx35600, nx35610, 
         nx35620, nx35630, nx35640, nx35650, nx35660, nx35670, nx35680, nx35690, 
         nx35700, nx35710, nx35720, nx35730, nx35740, nx35750, nx35760, nx35770, 
         nx35780, nx35790, nx35800, nx35810, nx35820, nx35830, nx35840, nx35850, 
         nx35860, nx35870, nx35880, nx35890, nx35900, nx35910, nx35920, nx35930, 
         nx35940, nx35950, nx35960, nx35970, nx35980, nx35990, nx36000, nx36010, 
         nx36020, nx36030, nx36040, nx36050, nx36060, nx36070, nx36080, nx36090, 
         nx36100, nx36110, nx36120, nx36130, nx36140, nx36150, nx36160, nx36170, 
         nx36180, nx36190, nx36200, nx36210, nx36220, nx36230, nx36240, nx36250, 
         nx36260, nx36270, nx36280, nx36290, nx36300, nx36310, nx36320, nx36330, 
         nx36340, nx36350, nx36360, nx36370, nx36380, nx36390, nx36400, nx36410, 
         nx36420, nx36430, nx36440, nx36450, nx36460, nx36470, nx36480, nx36490, 
         nx36500, nx36510, nx36520, nx36530, nx36540, nx36550, nx36560, nx36570, 
         nx36580, nx36590, nx36600, nx36610, nx36620, nx36630, nx36640, nx36650, 
         nx36660, nx36670, nx36680, nx36690, nx36700, nx36710, nx36720, nx36730, 
         nx36740, nx36750, nx36760, nx36770, nx36780, nx36790, nx36800, nx36810, 
         nx36820, nx36830, nx36840, nx36850, nx36860, nx36870, nx36880, nx36890, 
         nx36900, nx36910, nx36920, nx36930, nx36940, nx36950, nx36960, nx36970, 
         nx36980, nx36990, nx37000, nx37010, nx37020, nx37030, nx37040, nx37050, 
         nx37060, nx37070, nx37080, nx37090, nx37100, nx37110, nx37120, nx37130, 
         nx37140, nx37150, nx37160, nx37170, nx37180, nx37190, nx37200, nx37210, 
         nx37220, nx37230, nx37240, nx37250, nx37260, nx37270, nx37280, nx37290, 
         nx37300, nx37310, nx37320, nx37330, nx37340, nx37350, nx37360, nx37370, 
         nx37380, nx37390, nx37400, nx37410, nx37420, nx37430, nx37440, nx37450, 
         nx37460, nx37470, nx37480, nx37490, nx37500, nx37510, nx37520, nx37530, 
         nx37540, nx37550, nx37560, nx37570, nx37580, nx37590, nx37600, nx37610, 
         nx37620, nx37630, nx37640, nx37650, nx37660, nx37670, nx37680, nx37690, 
         nx37700, nx37710, nx37720, nx37730, nx37740, nx37750, nx37760, nx37770, 
         nx37780, nx37790, nx37800, nx37810, nx37820, nx37830, nx37840, nx37850, 
         nx37860, nx37870, nx37880, nx37890, nx37900, nx37910, nx37920, nx37930, 
         nx37940, nx37950, nx37960, nx37970, nx37980, nx37990, nx38000, nx38010, 
         nx38020, nx38030, nx38040, nx38050, nx38060, nx38070, nx38080, nx38090, 
         nx38100, nx38110, nx38120, nx38130, nx38140, nx38150, nx38160, nx38170, 
         nx38180, nx38190, nx38200, nx38210, nx38220, nx38230, nx38240, nx38250, 
         nx38260, nx38270, nx38280, nx38290, nx38300, nx38310, nx38320, nx38330, 
         nx38340, nx38350, nx38360, nx38370, nx38380, nx38390, nx38400, nx38410, 
         nx38420, nx38430, nx38440, nx38450, nx38460, nx38470, nx38480, nx38490, 
         nx38500, nx38510, nx38520, nx38530, nx38540, nx38550, nx38560, nx38570, 
         nx38580, nx38590, nx38600, nx38610, nx38620, nx38630, nx38640, nx38650, 
         nx38660, nx38670, nx38680, nx38690, nx38700, nx38710, nx38720, nx38730, 
         nx38740, nx38750, nx38760, nx38770, nx38780, nx38790, nx38800, nx38810, 
         nx38820, nx38830, nx38840, nx38850, nx38860, nx38870, nx38880, nx38890, 
         nx38900, nx38910, nx38920, nx38930, nx38940, nx38950, nx38960, nx38970, 
         nx38980, nx38990, nx39000, nx39010, nx39020, nx39030, nx39040, nx39050, 
         nx39060, nx39070, nx39080, nx39090, nx39100, nx39110, nx39120, nx39130, 
         nx39140, nx39150, nx39160, nx39170, nx39180, nx39190, nx39200, nx39210, 
         nx39220, nx39230, nx39240, nx39250, nx39260, nx39270, nx39280, nx39290, 
         nx39300, nx39310, nx39320, nx39330, nx39340, nx39350, nx39360, nx39370, 
         nx39380, nx39390, nx39400, nx39410, nx39420, nx39430, nx39440, nx39450, 
         nx39460, nx39470, nx39480, nx39490, nx39500, nx39510, nx39520, nx39530, 
         nx39540, nx39550, nx39560, nx39570, nx39580, nx39590, nx39600, nx39610, 
         nx39620, nx39630, nx39640, nx39650, nx39660, nx39670, nx39680, nx39690, 
         nx39700, nx39710, nx39720, nx39730, nx39740, nx39750, nx39760, nx39770, 
         nx39780, nx39790, nx39800, nx39810, nx39820, nx39830, nx39840, nx39850, 
         nx39860, nx39870, nx39880, nx39890, nx39900, nx39910, nx39920, nx39930, 
         nx39940, nx39950, nx39960, nx39970, nx39980, nx39990, nx40000, nx40010, 
         nx40020, nx40030, nx40040, nx40050, nx40060, nx40070, nx40080, nx40090, 
         nx40100, nx40110, nx40120, nx40130, nx40140, nx40150, nx40160, nx40170, 
         nx40180, nx40190, nx40200, nx40210, nx40220, nx40230, nx40240, nx40250, 
         nx40260, nx40270, nx40280, nx40290, nx40300, nx40310, nx40320, nx40330, 
         nx40340, nx40350, nx40360, nx40370, nx40380, nx40390, nx40400, nx40410, 
         nx40420, nx40430, nx40440, nx40450, nx40460, nx40470, nx40480, nx40490, 
         nx40500, nx40510, nx40520, nx40530, nx40540, nx40550, nx40560, nx40570, 
         nx40580, nx40590, nx40600, nx40610, nx40620, nx40630, nx40640, nx40650, 
         nx40660, nx40670, nx40680, nx40690, nx40700, nx40710, nx40720, nx40730, 
         nx40740, nx40750, nx40760, nx40770, nx40780, nx40790, nx40800, nx40810, 
         nx40820, nx40830, nx40840, nx40850, nx40860, nx40870, nx40880, nx40890, 
         nx40900, nx40910, nx40920, nx40930, nx40940, nx40950, nx40960, nx40970, 
         nx40980, nx40990, nx41000, nx41010, nx41020, nx41030, nx41040, nx41050, 
         nx41060, nx41070, nx41080, nx41090, nx41100, nx41110, nx41120, nx41130, 
         nx41140, nx41150, nx41160, nx41170, nx41180, nx41190, nx41200, nx41210, 
         nx41220, nx41230, nx41240, nx41250, nx41260, nx41270, nx41280, nx41290, 
         nx41300, nx41310, nx41320, nx41330, nx41340, nx41350, nx41360, nx41370, 
         nx41380, nx41390, nx41400, nx41410, nx41420, nx41430, nx41440, nx41450, 
         nx41460, nx41470, nx41480, nx41490, nx41500, nx41510, nx41520, nx41530, 
         nx41540, nx41550, nx41560, nx41570, nx41580, nx41590, nx41600, nx41610, 
         nx41620, nx41630, nx41640, nx41650, nx41660, nx41670, nx41680, nx41690, 
         nx41700, nx41710, nx41720, nx41730, nx41740, nx41750, nx41760, nx41770, 
         nx41780, nx41790, nx41800, nx41810, nx41820, nx41830, nx41840, nx41850, 
         nx41860, nx41870, nx41880, nx41890, nx41900, nx41910, nx41920, nx41930, 
         nx41940, nx41950, nx41960, nx41970, nx41980, nx41990, nx42000, nx42010, 
         nx42020, nx42030, nx42040, nx42050, nx42060, nx42070, nx42080, nx42090, 
         nx42100, nx42110, nx42120, nx42130, nx42140, nx42150, nx42160, nx42170, 
         nx42180, nx42190, nx42200, nx42210, nx42220, nx42230, nx42240, nx42250, 
         nx42260, nx42270, nx42280, nx42290, nx42300, nx42310, nx42320, nx42330, 
         nx42340, nx42350, nx42360, nx42370, nx42380, nx42390, nx42400, nx42410, 
         nx42420, nx42430, nx42440, nx42450, nx42460, nx42470, nx42480, nx42490, 
         nx42500, nx42510, nx42520, nx42530, nx42540, nx42550, nx42560, nx42570, 
         nx42580, nx42590, nx42600, nx42610, nx42620, nx42630, nx42640, nx42650, 
         nx42660, nx42670, nx42680, nx42690, nx42700, nx42710, nx42720, nx42730, 
         nx42740, nx42750, nx42760, nx42770, nx42780, nx42790, nx42800, nx42810, 
         nx42820, nx42830, nx42840, nx42850, nx42860, nx42870, nx42880, nx42890, 
         nx42900, nx42910, nx42920, nx42930, nx42940, nx42950, nx42960, nx42970, 
         nx42980, nx42990, nx43000, nx43010, nx43020, nx43030, nx43040, nx43050, 
         nx43060, nx43070, nx43080, nx43090, nx43100, nx43110, nx43120, nx43130, 
         nx43140, nx43150, nx43160, nx43170, nx43180, nx43190, nx43200, nx43210, 
         nx43220, nx43230, nx43240, nx43250, nx43260, nx43270, nx43280, nx43290, 
         nx43300, nx43310, nx43320, nx43330, nx43340, nx43350, nx43360, nx43370, 
         nx43380, nx43390, nx43400, nx43410, nx43420, nx43430, nx43440, nx43450, 
         nx43460, nx43470, nx43480, nx43490, nx43500, nx43510, nx43520, nx43530, 
         nx43540, nx43550, nx43560, nx43570, nx43580, nx43590, nx43600, nx43610, 
         nx43620, nx43630, nx43640, nx43650, nx43660, nx43670, nx43680, nx43690, 
         nx43700, nx43710, nx43720, nx43730, nx43740, nx43750, nx43760, nx43770, 
         nx43780, nx43790, nx43800, nx43810, nx43820, nx43830, nx43840, nx43850, 
         nx43860, nx43870, nx43880, nx43890, nx43900, nx43910, nx43920, nx43930, 
         nx43940, nx43950, nx43960, nx43970, nx43980, nx43990, nx44000, nx44010, 
         nx44020, nx44030, nx44040, nx44050, nx44060, nx44070, nx44080, nx44090, 
         nx44100, nx44110, nx44120, nx44130, nx44140, nx44150, nx44160, nx44170, 
         nx44180, nx44190, nx44200, nx44210, nx44220, nx44230, nx44240, nx44250, 
         nx44260, nx44270, nx44280, nx44290, nx44300, nx44310, nx44320, nx44330, 
         nx44340, nx44350, nx44360, nx44370, nx44380, nx44390, nx44400, nx44410, 
         nx44420, nx44430, nx44440, nx44450, nx44460, nx44470, nx44480, nx44490, 
         nx44500, nx44510, nx44520, nx44530, nx44540, nx44550, nx44560, nx44570, 
         nx44580, nx44590, nx44600, nx44610, nx44620, nx44630, nx44640, nx44650, 
         nx44660, nx44670, nx44680, nx44690, nx44700, nx44710, nx44720, nx44730, 
         nx44740, nx44750, nx44760, nx44770, nx44780, nx44790, nx44800, nx44810, 
         nx44820, nx44830, nx44840, nx44850, nx44860, nx44870, nx44880, nx44890, 
         nx44900, nx44910, nx44920, nx44930, nx44940, nx44950, nx44960, nx44970, 
         nx44980, nx44990, nx45000, nx45010, nx45020, nx45030, nx45040, nx45050, 
         nx45060, nx45070, nx45080, nx45090, nx45100, nx45110, nx45120, nx45130, 
         nx45140, nx45150, nx45160, nx45170, nx45180, nx45190, nx45200, nx45210, 
         nx45220, nx45230, nx45240, nx45250, nx45260, nx45270, nx45280, nx45290, 
         nx45300, nx45310, nx45320, nx45330, nx45340, nx45350, nx45360, nx45370, 
         nx45380, nx45390, nx45400, nx45410, nx45420, nx45430, nx45440, nx45450, 
         nx45460, nx45470, nx45480, nx45490, nx45500, nx45510, nx45520, nx45530, 
         nx45540, nx45550, nx45560, nx45570, nx45580, nx45590, nx45600, nx45610, 
         nx45620, nx45630, nx45640, nx45650, nx45660, nx45670, nx45680, nx45690, 
         nx45700, nx45710, nx45720, nx45730, nx45740, nx45750, nx45760, nx45770, 
         nx45780, nx45790, nx45800, nx45810, nx45820, nx45830, nx45840, nx45850, 
         nx45860, nx45870, nx45880, nx45890, nx45900, nx45910, nx45920, nx45930, 
         nx45940, nx45950, nx45960, nx45970, nx45980, nx45990, nx46000, nx46010, 
         nx46020, nx46030, nx46040, nx46050, nx46060, nx46070, nx46080, nx46090, 
         nx46100, nx46110, nx46120, nx46130, nx46140, nx46150, nx46160, nx46170, 
         nx46180, nx46190, nx46200, nx46210, nx46220, nx46230, nx46240, nx46250, 
         nx46260, nx46270, nx46280, nx46290, nx46300, nx46310, nx46320, nx46330, 
         nx46340, nx46350, nx46360, nx46370, nx46380, nx46390, nx46400, nx46410, 
         nx46420, nx46430, nx46440, nx46450, nx46460, nx46470, nx46480, nx46490, 
         nx46500, nx46510, nx46520, nx46530, nx46540, nx46550, nx46560, nx46570, 
         nx46580, nx46590, nx46600, nx46610, nx46620, nx46630, nx46640, nx46650, 
         nx46660, nx46670, nx46680, nx46690, nx46700, nx46710, nx46720, nx46730, 
         nx46740, nx46750, nx46760, nx46770, nx46780, nx46790, nx46800, nx46810, 
         nx46820, nx46830, nx46840, nx46850, nx46860, nx46870, nx46880, nx46890, 
         nx46900, nx46910, nx46920, nx46930, nx46940, nx46950, nx46960, nx46970, 
         nx46980, nx46990, nx47000, nx47010, nx47020, nx47030, nx47040, nx47050, 
         nx47060, nx47070, nx47080, nx47090, nx47100, nx47110, nx47120, nx47130, 
         nx47140, nx47150, nx47160, nx47170, nx47180, nx47190, nx47200, nx47210, 
         nx47220, nx47230, nx47240, nx47250, nx47260, nx47270, nx47280, nx47290, 
         nx47300, nx47310, nx47320, nx47330, nx47340, nx47350, nx47360, nx47370, 
         nx47380, nx47390, nx47400, nx47410, nx47420, nx47430, nx47440, nx47450, 
         nx47460, nx47470, nx47480, nx47490, nx47500, nx47510, nx47520, nx47530, 
         nx47540, nx47550, nx47560, nx47570, nx47580, nx47590, nx47600, nx47610, 
         nx47620, nx47630, nx47640, nx47650, nx47660, nx47670, nx47680, nx47690, 
         nx47700, nx47710, nx47720, nx47730, nx47740, nx47750, nx47760, nx47770, 
         nx47780, nx47790, nx47800, nx47810, nx47820, nx47830, nx47840, nx47850, 
         nx47860, nx47870, nx47880, nx47890, nx47900, nx47910, nx47920, nx47930, 
         nx47940, nx47950, nx47960, nx47970, nx47980, nx47990, nx48000, nx48010, 
         nx48020, nx48030, nx48040, nx48050, nx48060, nx48070, nx48080, nx48090, 
         nx48100, nx48110, nx48120, nx48130, nx48140, nx48150, nx48160, nx48170, 
         nx48180, nx48190, nx48200, nx48210, nx48220, nx48230, nx48240, nx48250, 
         nx48260, nx48270, nx48280, nx48290, nx48300, nx48310, nx48320, nx48330, 
         nx48340, nx48350, nx48360, nx48370, nx48380, nx48390, nx48400, nx48410, 
         nx48420, nx48430, nx48440, nx48450, nx48460, nx48470, nx48480, nx48490, 
         nx48500, nx48510, nx48520, nx48530, nx48540, nx48550, nx48560, nx48570, 
         nx48580, nx48590, nx48600, nx48610, nx48620, nx48630, nx48640, nx48650, 
         nx48660, nx48670, nx48680, nx48690, nx48700, nx48710, nx48720, nx48730, 
         nx48740, nx48750, nx48760, nx48770, nx48780, nx48790, nx48800, nx48810, 
         nx48820, nx48830, nx48840, nx48850, nx48860, nx48870, nx48880, nx48890, 
         nx48900, nx48910, nx48920, nx48930, nx48940, nx48950, nx48960, nx48970, 
         nx48980, nx48990, nx49000, nx49010, nx49020, nx49030, nx49040, nx49050, 
         nx49060, nx49070, nx49080, nx49090, nx49100, nx49110, nx49120, nx49130, 
         nx49140, nx49150, nx49160, nx49170, nx49180, nx49190, nx49200, nx49210, 
         nx49220, nx49230, nx49240, nx49250, nx49260, nx49270, nx49280, nx49290, 
         nx49300, nx49310, nx49320, nx49330, nx49340, nx49350, nx49360, nx49370, 
         nx49380, nx49390, nx49400, nx49410, nx49420, nx49430, nx49440, nx49450, 
         nx49460, nx49470, nx49480, nx49490, nx49500, nx49510, nx49520, nx49530, 
         nx49540, nx49550, nx49560, nx49570, nx49580, nx49590, nx49600, nx49610, 
         nx49620, nx49630, nx49640, nx49650, nx49660, nx49670, nx49680, nx49690, 
         nx49700, nx49710, nx49720, nx49730, nx49740, nx49750, nx49760, nx49770, 
         nx49780, nx49790, nx49800, nx49810, nx49820, nx49830, nx49840, nx49850, 
         nx49860, nx49870, nx49880, nx49890, nx49900, nx49910, nx49920, nx49930, 
         nx49940, nx49950, nx49960, nx49970, nx49980, nx49990, nx50000, nx50010, 
         nx50020, nx50030, nx50040, nx50050, nx50060, nx50070, nx50080, nx50090, 
         nx50100, nx50110, nx50120, nx50130, nx50140, nx50150, nx50160, nx50170, 
         nx50180, nx50190, nx50200, nx50210, nx50220, nx50230, nx50240, nx50250, 
         nx50260, nx50270, nx50280, nx50290, nx50300, nx50310, nx50320, nx50330, 
         nx50340, nx50350, nx50360, nx50370, nx50380, nx50390, nx50400, nx50410, 
         nx50420, nx50430, nx50440, nx50450, nx50460, nx50470, nx50480, nx50490, 
         nx50500, nx50510, nx50520, nx50530, nx50540, nx50550, nx50560, nx50570, 
         nx50580, nx50590, nx50600, nx50610, nx50620, nx50630, nx50640, nx50650, 
         nx50660, nx50670, nx50680, nx50690, nx50700, nx50710, nx50720, nx50730, 
         nx50740, nx50750, nx50760, nx50770, nx50780, nx50790, nx50800, nx50810, 
         nx50820, nx50830, nx50840, nx50850, nx50860, nx50870, nx50880, nx50890, 
         nx50900, nx50910, nx50920, nx50930, nx50940, nx50950, nx50960, nx50970, 
         nx50980, nx50990, nx51000, nx51010, nx51020, nx51030, nx51040, nx51050, 
         nx51060, nx51070, nx51080, nx51090, nx51100, nx51110, nx51120, nx51130, 
         nx51140, nx51150, nx51160, nx51170, nx51180, nx51190, nx51200, nx51210, 
         nx51220, nx51230, nx51240, nx51250, nx51260, nx51270, nx51280, nx51290, 
         nx51300, nx51310, nx51320, nx51330, nx51340, nx51350, nx51360, nx51370, 
         nx51380, nx51390, nx51400, nx51410, nx51420, nx51430, nx51440, nx51450, 
         nx51460, nx51470, nx51480, nx51490, nx51500, nx51510, nx51520, nx51530, 
         nx51540, nx51550, nx51560, nx51570, nx51580, nx51590, nx51600, nx51610, 
         nx51620, nx51630, nx51640, nx51650, nx51660, nx51670, nx51680, nx51690, 
         nx51700, nx51710, nx51720, nx51730, nx51740, nx51750, nx51760, nx51770, 
         nx51780, nx51790, nx51800, nx51810, nx51820, nx51830, nx51840, nx51850, 
         nx51860, nx51870, nx51880, nx51890, nx51900, nx51910, nx51920, nx51930, 
         nx51940, nx51950, nx51960, nx51970, nx51980, nx51990, nx52000, nx52010, 
         nx52020, nx52030, nx52040, nx52050, nx52060, nx52070, nx52080, nx52090, 
         nx52100, nx52110, nx52120, nx52130, nx52140, nx52150, nx52160, nx52170, 
         nx52180, nx52190, nx52200, nx52210, nx52220, nx52230, nx52240, nx52250, 
         nx52260, nx52270, nx52280, nx52290, nx52300, nx52310, nx52320, nx52330, 
         nx52340, nx52350, nx52360, nx52370, nx52380, nx52390, nx52400, nx52410, 
         nx52420, nx52430, nx52440, nx52450, nx52460, nx52470, nx52480, nx52490, 
         nx52500, nx52510, nx52520, nx52530, nx52540, nx52550, nx52560, nx52570, 
         nx52580, nx52590, nx52600, nx52610, nx52620, nx52630, nx52640, nx52650, 
         nx52660, nx52670, nx52680, nx52690, nx52700, nx52710, nx52720, nx52730, 
         nx52740, nx52750, nx52760, nx52770, nx52780, nx52790, nx52800, nx52810, 
         nx52820, nx52830, nx52840, nx52850, nx52860, nx52870, nx52880, nx52890, 
         nx52900, nx52910, nx52920, nx52930, nx52940, nx52950, nx52960, nx52970, 
         nx52980, nx52990, nx53000, nx53010, nx53020, nx53030, nx53040, nx53050, 
         nx53060, nx53070, nx53080, nx53090, nx53100, nx53110, nx53120, nx53130, 
         nx53140, nx53150, nx53160, nx53170, nx53180, nx53190, nx53200, nx53210, 
         nx53220, nx53230, nx53240, nx53250, nx53260, nx53270, nx53280, nx53290, 
         nx53300, nx53310, nx53320, nx53330, nx53340, nx53350, nx53360, nx53370, 
         nx53380, nx53390, nx53400, nx53410, nx53420, nx53430, nx53440, nx53450, 
         nx53460, nx53470, nx53480, nx53490, nx53500, nx53510, nx53520, nx53530, 
         nx53540, nx53550, nx53560, nx53570, nx53580, nx53590, nx53600, nx53610, 
         nx53620, nx53630, nx53640, nx53650, nx53660, nx53670, nx53680, nx53690, 
         nx53700, nx53710, nx53720, nx53730, nx53740, nx53750, nx53760, nx53770, 
         nx53780, nx53790, nx53800, nx53810, nx53820, nx53830, nx53840, nx53850, 
         nx53860, nx53870, nx53880, nx53890, nx53900, nx53910, nx53920, nx53930, 
         nx53940, nx53950, nx53960, nx53970, nx53980, nx53990, nx54000, nx54010, 
         nx54020, nx54030, nx54040, nx54050, nx54060, nx54070, nx54080, nx54090, 
         nx54100, nx54112, nx54115, nx54124, nx54126, nx54129, nx54135, nx54142, 
         nx54156, nx54163, nx54169, nx54183, nx54200, nx54206, nx54220, nx54236, 
         nx54253, nx54273, nx54276, nx54282, nx54291, nx54301, nx54311, nx54322, 
         nx54332, nx54342, nx54352, nx54364, nx54367, nx54373, nx54382, nx54392, 
         nx54402, nx54413, nx54423, nx54433, nx54443, nx54455, nx54458, nx54464, 
         nx54471, nx54481, nx54491, nx54502, nx54512, nx54522, nx54532, nx54545, 
         nx54548, nx54554, nx54563, nx54573, nx54583, nx54594, nx54604, nx54614, 
         nx54624, nx54636, nx54639, nx54650, nx54660, nx54670, nx54681, nx54691, 
         nx54701, nx54711, nx54723, nx54726, nx54732, nx54739, nx54749, nx54759, 
         nx54770, nx54780, nx54790, nx54800, nx54812, nx54815, nx54826, nx54836, 
         nx54846, nx54857, nx54867, nx54877, nx54887, nx54900, nx54903, nx54914, 
         nx54924, nx54934, nx54945, nx54955, nx54965, nx54975, nx54987, nx54990, 
         nx54994, nx54996, nx55001, nx55004, nx55008, nx55013, nx55016, nx55020, 
         nx55025, nx55028, nx55032, nx55037, nx55041, nx55045, nx55050, nx55053, 
         nx55057, nx55062, nx55065, nx55069, nx55074, nx55077, nx55081, nx55086, 
         nx55089, nx55092, nx55103, nx55113, nx55123, nx55134, nx55144, nx55154, 
         nx55164, nx55176, nx55179, nx55190, nx55200, nx55210, nx55221, nx55231, 
         nx55241, nx55251, nx55264, nx55267, nx55273, nx55282, nx55292, nx55302, 
         nx55313, nx55323, nx55333, nx55343, nx55355, nx55358, nx55369, nx55379, 
         nx55389, nx55400, nx55410, nx55420, nx55430, nx55442, nx55445, nx55456, 
         nx55466, nx55476, nx55487, nx55497, nx55507, nx55517, nx55529, nx55532, 
         nx55543, nx55553, nx55563, nx55574, nx55584, nx55594, nx55604, nx55618, 
         nx55621, nx55629, nx55637, nx55645, nx55654, nx55662, nx55670, nx55678, 
         nx55686, nx55689, nx55697, nx55705, nx55713, nx55722, nx55730, nx55738, 
         nx55746, nx55754, nx55757, nx55765, nx55773, nx55781, nx55790, nx55798, 
         nx55806, nx55814, nx55822, nx55825, nx55833, nx55841, nx55849, nx55858, 
         nx55866, nx55874, nx55882, nx55891, nx55894, nx55902, nx55910, nx55918, 
         nx55927, nx55935, nx55943, nx55951, nx55959, nx55962, nx55970, nx55978, 
         nx55986, nx55995, nx56003, nx56011, nx56019, nx56027, nx56030, nx56038, 
         nx56046, nx56054, nx56063, nx56071, nx56079, nx56087, nx56095, nx56098, 
         nx56106, nx56114, nx56122, nx56131, nx56139, nx56147, nx56155, nx56164, 
         nx56167, nx56175, nx56183, nx56191, nx56200, nx56208, nx56216, nx56224, 
         nx56232, nx56235, nx56243, nx56251, nx56259, nx56268, nx56276, nx56284, 
         nx56292, nx56300, nx56303, nx56311, nx56319, nx56327, nx56336, nx56344, 
         nx56352, nx56360, nx56368, nx56371, nx56379, nx56387, nx56395, nx56404, 
         nx56412, nx56420, nx56428, nx56437, nx56440, nx56448, nx56456, nx56464, 
         nx56473, nx56481, nx56489, nx56497, nx56505, nx56508, nx56516, nx56524, 
         nx56532, nx56541, nx56549, nx56557, nx56565, nx56573, nx56576, nx56584, 
         nx56592, nx56600, nx56609, nx56617, nx56625, nx56633, nx56641, nx56644, 
         nx56652, nx56660, nx56668, nx56677, nx56685, nx56693, nx56701, nx56711, 
         nx56714, nx56722, nx56730, nx56738, nx56747, nx56755, nx56763, nx56771, 
         nx56779, nx56782, nx56790, nx56798, nx56806, nx56815, nx56823, nx56831, 
         nx56839, nx56847, nx56850, nx56858, nx56866, nx56874, nx56883, nx56891, 
         nx56899, nx56907, nx56915, nx56918, nx56926, nx56934, nx56942, nx56951, 
         nx56959, nx56967, nx56975, nx56984, nx56987, nx56995, nx57003, nx57011, 
         nx57020, nx57028, nx57036, nx57044, nx57052, nx57055, nx57063, nx57071, 
         nx57079, nx57088, nx57096, nx57104, nx57112, nx57120, nx57123, nx57131, 
         nx57139, nx57147, nx57156, nx57164, nx57172, nx57180, nx57188, nx57191, 
         nx57199, nx57207, nx57215, nx57224, nx57232, nx57240, nx57248, nx57257, 
         nx57260, nx57268, nx57276, nx57284, nx57293, nx57301, nx57309, nx57317, 
         nx57325, nx57328, nx57336, nx57344, nx57352, nx57361, nx57369, nx57377, 
         nx57385, nx57393, nx57396, nx57404, nx57412, nx57420, nx57429, nx57437, 
         nx57445, nx57453, nx57461, nx57464, nx57472, nx57480, nx57488, nx57497, 
         nx57505, nx57513, nx57521, nx57530, nx57533, nx57541, nx57549, nx57557, 
         nx57566, nx57574, nx57582, nx57590, nx57598, nx57601, nx57609, nx57617, 
         nx57625, nx57634, nx57642, nx57650, nx57658, nx57666, nx57669, nx57677, 
         nx57685, nx57693, nx57702, nx57710, nx57718, nx57726, nx57734, nx57737, 
         nx57745, nx57753, nx57761, nx57770, nx57778, nx57786, nx57794, nx57804, 
         nx57807, nx57815, nx57823, nx57831, nx57840, nx57848, nx57856, nx57864, 
         nx57872, nx57875, nx57883, nx57891, nx57899, nx57908, nx57916, nx57924, 
         nx57932, nx57940, nx57943, nx57951, nx57959, nx57967, nx57976, nx57984, 
         nx57992, nx58000, nx58008, nx58011, nx58019, nx58027, nx58035, nx58044, 
         nx58052, nx58060, nx58068, nx58077, nx58080, nx58088, nx58096, nx58104, 
         nx58113, nx58121, nx58129, nx58137, nx58145, nx58148, nx58156, nx58164, 
         nx58172, nx58181, nx58189, nx58197, nx58205, nx58213, nx58216, nx58224, 
         nx58232, nx58240, nx58249, nx58257, nx58265, nx58273, nx58281, nx58284, 
         nx58292, nx58300, nx58308, nx58317, nx58325, nx58333, nx58341, nx58350, 
         nx58353, nx58361, nx58369, nx58377, nx58386, nx58394, nx58402, nx58410, 
         nx58418, nx58421, nx58429, nx58437, nx58445, nx58454, nx58462, nx58470, 
         nx58478, nx58486, nx58489, nx58497, nx58505, nx58513, nx58522, nx58530, 
         nx58538, nx58546, nx58554, nx58557, nx58565, nx58573, nx58581, nx58590, 
         nx58598, nx58606, nx58614, nx58623, nx58626, nx58634, nx58642, nx58650, 
         nx58659, nx58667, nx58675, nx58683, nx58691, nx58694, nx58702, nx58710, 
         nx58718, nx58727, nx58735, nx58743, nx58751, nx58759, nx58762, nx58770, 
         nx58778, nx58786, nx58795, nx58803, nx58811, nx58819, nx58827, nx58830, 
         nx58838, nx58846, nx58854, nx58863, nx58871, nx58879, nx58887, nx58897, 
         nx58900, nx58908, nx58916, nx58924, nx58933, nx58941, nx58949, nx58957, 
         nx58965, nx58968, nx58976, nx58984, nx58992, nx59001, nx59009, nx59017, 
         nx59025, nx59033, nx59036, nx59044, nx59052, nx59060, nx59069, nx59077, 
         nx59085, nx59093, nx59101, nx59104, nx59112, nx59120, nx59128, nx59137, 
         nx59145, nx59153, nx59161, nx59170, nx59173, nx59181, nx59189, nx59197, 
         nx59206, nx59214, nx59222, nx59230, nx59238, nx59241, nx59249, nx59257, 
         nx59265, nx59274, nx59282, nx59290, nx59298, nx59306, nx59309, nx59317, 
         nx59325, nx59333, nx59342, nx59350, nx59358, nx59366, nx59374, nx59377, 
         nx59385, nx59393, nx59401, nx59410, nx59418, nx59426, nx59434, nx59443, 
         nx59446, nx59454, nx59462, nx59470, nx59479, nx59487, nx59495, nx59503, 
         nx59511, nx59514, nx59522, nx59530, nx59538, nx59547, nx59555, nx59563, 
         nx59571, nx59579, nx59582, nx59590, nx59598, nx59606, nx59615, nx59623, 
         nx59631, nx59639, nx59647, nx59650, nx59658, nx59666, nx59674, nx59683, 
         nx59691, nx59699, nx59707, nx59716, nx59719, nx59727, nx59735, nx59743, 
         nx59752, nx59760, nx59768, nx59776, nx59784, nx59787, nx59795, nx59803, 
         nx59811, nx59820, nx59828, nx59836, nx59844, nx59852, nx59855, nx59863, 
         nx59871, nx59879, nx59888, nx59896, nx59904, nx59912, nx59920, nx59923, 
         nx59931, nx59939, nx59947, nx59956, nx59964, nx59972, nx59980, nx59990, 
         nx59993, nx60001, nx60009, nx60017, nx60026, nx60034, nx60042, nx60050, 
         nx60058, nx60061, nx60069, nx60077, nx60085, nx60094, nx60102, nx60110, 
         nx60118, nx60126, nx60129, nx60137, nx60145, nx60153, nx60162, nx60170, 
         nx60178, nx60186, nx60194, nx60197, nx60205, nx60213, nx60221, nx60230, 
         nx60238, nx60246, nx60254, nx60263, nx60266, nx60274, nx60282, nx60290, 
         nx60299, nx60307, nx60315, nx60323, nx60331, nx60334, nx60342, nx60350, 
         nx60358, nx60367, nx60375, nx60383, nx60391, nx60399, nx60402, nx60410, 
         nx60418, nx60426, nx60435, nx60443, nx60451, nx60459, nx60467, nx60470, 
         nx60478, nx60486, nx60494, nx60503, nx60511, nx60519, nx60527, nx60536, 
         nx60539, nx60547, nx60555, nx60563, nx60572, nx60580, nx60588, nx60596, 
         nx60604, nx60607, nx60615, nx60623, nx60631, nx60640, nx60648, nx60656, 
         nx60664, nx60672, nx60675, nx60683, nx60691, nx60699, nx60708, nx60716, 
         nx60724, nx60732, nx60740, nx60743, nx60751, nx60759, nx60767, nx60776, 
         nx60784, nx60792, nx60800, nx60809, nx60812, nx60820, nx60828, nx60836, 
         nx60845, nx60853, nx60861, nx60869, nx60877, nx60880, nx60888, nx60896, 
         nx60904, nx60913, nx60921, nx60929, nx60937, nx60945, nx60948, nx60956, 
         nx60964, nx60972, nx60981, nx60989, nx60997, nx61005, nx61013, nx61016, 
         nx61024, nx61032, nx61040, nx61049, nx61057, nx61065, nx61073, nx61083, 
         nx61086, nx61094, nx61102, nx61110, nx61119, nx61127, nx61135, nx61143, 
         nx61151, nx61154, nx61162, nx61170, nx61178, nx61187, nx61195, nx61203, 
         nx61211, nx61219, nx61222, nx61230, nx61238, nx61246, nx61255, nx61263, 
         nx61271, nx61279, nx61287, nx61290, nx61298, nx61306, nx61314, nx61323, 
         nx61331, nx61339, nx61347, nx61356, nx61359, nx61367, nx61375, nx61383, 
         nx61392, nx61400, nx61408, nx61416, nx61424, nx61427, nx61435, nx61443, 
         nx61451, nx61460, nx61468, nx61476, nx61484, nx61492, nx61495, nx61503, 
         nx61511, nx61519, nx61528, nx61536, nx61544, nx61552, nx61560, nx61563, 
         nx61571, nx61579, nx61587, nx61596, nx61604, nx61612, nx61620, nx61629, 
         nx61632, nx61640, nx61648, nx61656, nx61665, nx61673, nx61681, nx61689, 
         nx61697, nx61700, nx61708, nx61716, nx61724, nx61733, nx61741, nx61749, 
         nx61757, nx61765, nx61768, nx61776, nx61784, nx61792, nx61801, nx61809, 
         nx61817, nx61825, nx61833, nx61836, nx61844, nx61852, nx61860, nx61869, 
         nx61877, nx61885, nx61893, nx61902, nx61905, nx61913, nx61921, nx61929, 
         nx61938, nx61946, nx61954, nx61962, nx61970, nx61973, nx61981, nx61989, 
         nx61997, nx62006, nx62014, nx62022, nx62030, nx62038, nx62041, nx62049, 
         nx62057, nx62065, nx62074, nx62082, nx62090, nx62098, nx62106, nx62109, 
         nx62117, nx62125, nx62133, nx62142, nx62150, nx62158, nx62166, nx62176, 
         nx62179, nx62187, nx62195, nx62203, nx62212, nx62220, nx62228, nx62236, 
         nx62244, nx62247, nx62255, nx62263, nx62271, nx62280, nx62288, nx62296, 
         nx62304, nx62312, nx62315, nx62323, nx62331, nx62339, nx62348, nx62356, 
         nx62364, nx62372, nx62380, nx62383, nx62391, nx62399, nx62407, nx62416, 
         nx62424, nx62432, nx62440, nx62449, nx62452, nx62460, nx62468, nx62476, 
         nx62485, nx62493, nx62501, nx62509, nx62517, nx62520, nx62528, nx62536, 
         nx62544, nx62553, nx62561, nx62569, nx62577, nx62585, nx62588, nx62596, 
         nx62604, nx62612, nx62621, nx62629, nx62637, nx62645, nx62653, nx62656, 
         nx62664, nx62672, nx62680, nx62689, nx62697, nx62705, nx62713, nx62722, 
         nx62725, nx62733, nx62741, nx62749, nx62758, nx62766, nx62774, nx62782, 
         nx62790, nx62793, nx62801, nx62809, nx62817, nx62826, nx62834, nx62842, 
         nx62850, nx62858, nx62861, nx62869, nx62877, nx62885, nx62894, nx62902, 
         nx62910, nx62918, nx62926, nx62929, nx62937, nx62945, nx62953, nx62962, 
         nx62970, nx62978, nx62986, nx62995, nx62998, nx63006, nx63014, nx63022, 
         nx63031, nx63039, nx63047, nx63055, nx63063, nx63066, nx63074, nx63082, 
         nx63090, nx63099, nx63107, nx63115, nx63123, nx63131, nx63134, nx63142, 
         nx63150, nx63158, nx63167, nx63175, nx63183, nx63191, nx63199, nx63202, 
         nx63210, nx63218, nx63226, nx63235, nx63243, nx63251, nx63259, nx63284, 
         nx63286, nx63294, nx63296, nx63304, nx63306, nx63314, nx63316, nx63324, 
         nx63326, nx63334, nx63336, nx63344, nx63346, nx63354, nx63356, nx63364, 
         nx63366, nx63374, nx63376, nx63384, nx63386, nx63394, nx63396, nx63404, 
         nx63406, nx63414, nx63416, nx63424, nx63426, nx63434, nx63436, nx63444, 
         nx63446, nx63448, nx63450, nx63452, nx63454, nx63456, nx63458, nx63460, 
         nx63462, nx63464, nx63466, nx63468, nx63470, nx63472, nx63474, nx63476, 
         nx63478, nx63480, nx63482, nx63484, nx63486, nx63488, nx63490, nx63492, 
         nx63494, nx63496, nx63498, nx63500, nx63502, nx63504, nx63506, nx63514, 
         nx63516, nx63518, nx63520, nx63522, nx63524, nx63526, nx63528, nx63530, 
         nx63532, nx63534, nx63536, nx63538, nx63540, nx63542, nx63544, nx63546, 
         nx63548, nx63550, nx63552, nx63554, nx63556, nx63558, nx63560, nx63562, 
         nx63564, nx63566, nx63568, nx63570, nx63572, nx63574, nx63576, nx63584, 
         nx63586, nx63588, nx63590, nx63592, nx63594, nx63596, nx63598, nx63600, 
         nx63602, nx63604, nx63606, nx63608, nx63610, nx63612, nx63614, nx63616, 
         nx63618, nx63620, nx63622, nx63624, nx63626, nx63628, nx63630, nx63632, 
         nx63634, nx63636, nx63638, nx63640, nx63642, nx63644, nx63646, nx63654, 
         nx63656, nx63658, nx63660, nx63662, nx63664, nx63666, nx63668, nx63670, 
         nx63672, nx63674, nx63676, nx63678, nx63680, nx63682, nx63684, nx63686, 
         nx63688, nx63690, nx63692, nx63694, nx63696, nx63698, nx63700, nx63702, 
         nx63704, nx63706, nx63708, nx63710, nx63712, nx63714, nx63716, nx63724, 
         nx63726, nx63728, nx63730, nx63732, nx63734, nx63736, nx63738, nx63740, 
         nx63742, nx63744, nx63746, nx63748, nx63750, nx63752, nx63754, nx63756, 
         nx63758, nx63760, nx63762, nx63764, nx63766, nx63768, nx63770, nx63772, 
         nx63774, nx63776, nx63778, nx63780, nx63782, nx63784, nx63786, nx63794, 
         nx63796, nx63798, nx63800, nx63802, nx63804, nx63806, nx63808, nx63810, 
         nx63812, nx63814, nx63816, nx63818, nx63820, nx63822, nx63824, nx63826, 
         nx63828, nx63830, nx63832, nx63834, nx63836, nx63838, nx63840, nx63842, 
         nx63844, nx63846, nx63848, nx63850, nx63852, nx63854, nx63856, nx63864, 
         nx63866, nx63868, nx63870, nx63872, nx63874, nx63876, nx63878, nx63880, 
         nx63882, nx63884, nx63886, nx63888, nx63890, nx63892, nx63894, nx63896, 
         nx63898, nx63900, nx63902, nx63904, nx63906, nx63908, nx63910, nx63912, 
         nx63914, nx63916, nx63918, nx63920, nx63922, nx63924, nx63926, nx63934, 
         nx63936, nx63938, nx63940, nx63942, nx63944, nx63946, nx63948, nx63950, 
         nx63952, nx63954, nx63956, nx63958, nx63960, nx63962, nx63964, nx63966, 
         nx63968, nx63970, nx63972, nx63974, nx63976, nx63978, nx63980, nx63982, 
         nx63984, nx63986, nx63988, nx63990, nx63992, nx63994, nx63996, nx64004, 
         nx64006, nx64008, nx64010, nx64012, nx64014, nx64016, nx64018, nx64020, 
         nx64022, nx64024, nx64026, nx64028, nx64030, nx64032, nx64034, nx64036, 
         nx64038, nx64040, nx64042, nx64044, nx64046, nx64048, nx64050, nx64052, 
         nx64054, nx64056, nx64058, nx64060, nx64062, nx64064, nx64066, nx64074, 
         nx64076, nx64078, nx64080, nx64082, nx64084, nx64086, nx64088, nx64090, 
         nx64092, nx64094, nx64096, nx64098, nx64100, nx64102, nx64104, nx64106, 
         nx64108, nx64110, nx64112, nx64114, nx64116, nx64118, nx64120, nx64122, 
         nx64124, nx64126, nx64128, nx64130, nx64132, nx64134, nx64136, nx64144, 
         nx64146, nx64148, nx64150, nx64152, nx64154, nx64156, nx64158, nx64160, 
         nx64162, nx64164, nx64166, nx64168, nx64170, nx64172, nx64174, nx64176, 
         nx64178, nx64180, nx64182, nx64184, nx64186, nx64188, nx64190, nx64192, 
         nx64194, nx64196, nx64198, nx64200, nx64202, nx64204, nx64206, nx64214, 
         nx64216, nx64218, nx64220, nx64222, nx64224, nx64226, nx64228, nx64230, 
         nx64232, nx64234, nx64236, nx64238, nx64240, nx64242, nx64244, nx64246, 
         nx64248, nx64250, nx64252, nx64254, nx64256, nx64258, nx64260, nx64262, 
         nx64264, nx64266, nx64268, nx64270, nx64272, nx64274, nx64276, nx64284, 
         nx64286, nx64288, nx64290, nx64292, nx64294, nx64296, nx64298, nx64300, 
         nx64302, nx64304, nx64306, nx64308, nx64310, nx64312, nx64314, nx64316, 
         nx64318, nx64320, nx64322, nx64324, nx64326, nx64328, nx64330, nx64332, 
         nx64334, nx64336, nx64338, nx64340, nx64342, nx64344, nx64346, nx64354, 
         nx64356, nx64358, nx64360, nx64362, nx64364, nx64366, nx64368, nx64370, 
         nx64372, nx64374, nx64376, nx64378, nx64380, nx64382, nx64384, nx64386, 
         nx64388, nx64390, nx64392, nx64394, nx64396, nx64398, nx64400, nx64402, 
         nx64404, nx64406, nx64408, nx64410, nx64412, nx64414, nx64416, nx64488, 
         nx64490, nx64492, nx64494, nx64496, nx64498, nx64500, nx64502, nx64504, 
         nx64506, nx64508, nx64510, nx64512, nx64514, nx64516, nx64518, nx64520, 
         nx64522, nx64524, nx64526, nx64528, nx64530, nx64532, nx64534, nx64536, 
         nx64538, nx64540, nx64542, nx64544, nx64546, nx64548, nx64550, nx64552, 
         nx64554, nx64556, nx64558, nx64560, nx64562, nx64564, nx64566, nx64568, 
         nx64570, nx64572, nx64574, nx64576, nx64578, nx64580, nx64582, nx64584, 
         nx64586, nx64588, nx64590, nx64592, nx64594, nx64596, nx64598, nx64600, 
         nx64602, nx64604, nx64606, nx64608, nx64610, nx64612, nx64614, nx64616, 
         nx64618, nx64620, nx64622, nx64624, nx64626, nx64628, nx64630, nx64632, 
         nx64634, nx64636, nx64638, nx64640, nx64642, nx64644, nx64646, nx64648, 
         nx64650, nx64652, nx64654, nx64656, nx64658, nx64660, nx64662, nx64664, 
         nx64666, nx64668, nx64670, nx64672, nx64674, nx64676, nx64678, nx64680, 
         nx64682, nx64684, nx64686, nx64688, nx64690, nx64692, nx64694, nx64696, 
         nx64698, nx64700, nx64702, nx64704, nx64706, nx64708, nx64710, nx64712, 
         nx64714, nx64716, nx64718, nx64720, nx64722, nx64724, nx64726, nx64728, 
         nx64730, nx64732, nx64734, nx64736, nx64738, nx64740, nx64742, nx64744, 
         nx64746, nx64748, nx64750, nx64752, nx64754, nx64756, nx64758, nx64760, 
         nx64762, nx64764, nx64766, nx64768, nx64770, nx64772, nx64774, nx64776, 
         nx64778, nx64780, nx64782, nx64784, nx64786, nx64788, nx64790, nx64792, 
         nx64794, nx64796, nx64798, nx64800, nx64802, nx64804, nx64806, nx64808, 
         nx64810, nx64812, nx64814, nx64816, nx64818, nx64820, nx64822, nx64824, 
         nx64826, nx64828, nx64830, nx64832, nx64834, nx64836, nx64838, nx64840, 
         nx64842, nx64844, nx64846, nx64848, nx64850, nx64852, nx64854, nx64856, 
         nx64858, nx64860, nx64862, nx64864, nx64866, nx64868, nx64870, nx64872, 
         nx64874, nx64876, nx64878, nx64880, nx64882, nx64884, nx64886, nx64888, 
         nx64890, nx64892, nx64894, nx64896, nx64898, nx64900, nx64902, nx64904, 
         nx64906, nx64908, nx64910, nx64912, nx64914, nx64916, nx64918, nx64920, 
         nx64922, nx64924, nx64926, nx64928, nx64930, nx64932, nx64934, nx64936, 
         nx64938, nx64940, nx64942, nx64944, nx64946, nx64948, nx64950, nx64952, 
         nx64954, nx64956, nx64958, nx64960, nx64962, nx64964, nx64966, nx64968, 
         nx64970, nx64972, nx64974, nx64976, nx64978, nx64980, nx64982, nx64984, 
         nx64986, nx64988, nx64990, nx64992, nx64994, nx64996, nx64998, nx65000, 
         nx65002, nx65004, nx65006, nx65008, nx65010, nx65012, nx65014, nx65016, 
         nx65018, nx65020, nx65022, nx65024, nx65026, nx65028, nx65030, nx65032, 
         nx65034, nx65036, nx65038, nx65040, nx65042, nx65044, nx65046, nx65048, 
         nx65050, nx65052, nx65054, nx65056, nx65058, nx65060, nx65062, nx65064, 
         nx65066, nx65068, nx65070, nx65072, nx65074, nx65076, nx65078, nx65080, 
         nx65082, nx65084, nx65086, nx65088, nx65090, nx65092, nx65094, nx65096, 
         nx65098, nx65100, nx65102, nx65104, nx65106, nx65108, nx65110, nx65112, 
         nx65114, nx65116, nx65118, nx65120, nx65122, nx65124, nx65126, nx65128, 
         nx65130, nx65132, nx65134, nx65136, nx65138, nx65140, nx65142, nx65144, 
         nx65146, nx65148, nx65150, nx65152, nx65154, nx65156, nx65158, nx65160, 
         nx65162, nx65164, nx65166, nx65168, nx65170, nx65172, nx65174, nx65176, 
         nx65178, nx65180, nx65182, nx65184, nx65186, nx65188, nx65190, nx65192, 
         nx65194, nx65196, nx65198, nx65200, nx65202, nx65204, nx65206, nx65208, 
         nx65210, nx65212, nx65214, nx65216, nx65218, nx65220, nx65222, nx65224, 
         nx65226, nx65228, nx65234, nx65236, nx65238, nx65240, nx65242, nx65244, 
         nx65246, nx65248, nx65250, nx65252, nx65254, nx65256, nx65258, nx65260, 
         nx65262, nx65264, nx65266, nx65268, nx65270, nx65272, nx65274, nx65276, 
         nx65278, nx65280, nx65282, nx65284, nx65286, nx65288, nx65290, nx65292, 
         nx65294, nx65296, nx65298, nx65300, nx65302, nx65304, nx65306, nx65308, 
         nx65310, nx65312, nx65314, nx65316, nx65318, nx65320, nx65322, nx65324, 
         nx65326, nx65328, nx65330, nx65332, nx65334, nx65336, nx65338, nx65340, 
         nx65342, nx65344, nx65346, nx65348, nx65350, nx65352, nx65354, nx65356, 
         nx65358, nx65366, nx65368, nx65370, nx65372, nx65374, nx65376, nx65378, 
         nx65380, nx65382, nx65384, nx65386, nx65388, nx65390, nx65392, nx65394, 
         nx65396, nx65398, nx65400, nx65402, nx65404, nx65406, nx65408, nx65410, 
         nx65412, nx65414, nx65416, nx65418, nx65420, nx65422, nx65424, nx65426, 
         nx65428, nx65430, nx65432, nx65434, nx65436, nx65438, nx65440, nx65442, 
         nx65444, nx65446, nx65450, nx65452, nx65454, nx65456, nx65458, nx65460, 
         nx65462, nx65464, nx65466, nx65468, nx65470, nx65472, nx65474, nx65476, 
         nx65478, nx65480, nx65482, nx65484, nx65486, nx65488, nx65490, nx65492, 
         nx65494, nx65496, nx65498, nx65500, nx65502, nx65504, nx65506, nx65508, 
         nx65510, nx65512, nx65514, nx65516, nx65518, nx65520, nx65522, nx65526, 
         nx65528, nx65530, nx65532, nx65534, nx65536, nx65538, nx65540, nx65542, 
         nx65544, nx65546, nx65548, nx65550, nx65552, nx65554, nx65556, nx65558, 
         nx65560, nx65562, nx65564, nx65566, nx65568, nx65570, nx65572, nx65574, 
         nx65576, nx65578, nx65580, nx65582, nx65584, nx65586, nx65588, nx65590, 
         nx65592, nx65594, nx65596, nx65598, nx65602, nx65604, nx65606, nx65608, 
         nx65610, nx65612, nx65614, nx65616, nx65618, nx65620, nx65622, nx65624, 
         nx65626, nx65628, nx65630, nx65632, nx65634, nx65636, nx65638, nx65640, 
         nx65642, nx65644, nx65646, nx65648, nx65650, nx65652, nx65654, nx65656, 
         nx65658, nx65660, nx65662, nx65664, nx65666, nx65668, nx65670, nx65672, 
         nx65674, nx65678, nx65680, nx65682, nx65684, nx65686, nx65688, nx65690, 
         nx65692, nx65694, nx65696, nx65698, nx65700, nx65702, nx65704, nx65706, 
         nx65708, nx65710, nx65712, nx65714, nx65716, nx65718, nx65720, nx65722, 
         nx65724, nx65726, nx65728, nx65730, nx65732, nx65734, nx65736, nx65738, 
         nx65740, nx65742, nx65744, nx65746, nx65748, nx65750, nx65754, nx65756, 
         nx65758, nx65760, nx65762, nx65764, nx65766, nx65768, nx65770, nx65772, 
         nx65774, nx65776, nx65778, nx65780, nx65782, nx65784, nx65786, nx65788, 
         nx65790, nx65792, nx65794, nx65796, nx65798, nx65800, nx65802, nx65804, 
         nx65806, nx65808, nx65810, nx65812, nx65814, nx65816, nx65818, nx65820, 
         nx65822, nx65824, nx65826, nx65830, nx65832, nx65834, nx65836, nx65838, 
         nx65840, nx65842, nx65844, nx65846, nx65848, nx65850, nx65852, nx65854, 
         nx65856, nx65858, nx65860, nx65862, nx65864, nx65866, nx65868, nx65870, 
         nx65872, nx65874, nx65876, nx65878, nx65880, nx65882, nx65884, nx65886, 
         nx65888, nx65890, nx65892, nx65894, nx65896, nx65898, nx65900, nx65902, 
         nx65906, nx65908, nx65910, nx65912, nx65914, nx65916, nx65918, nx65920, 
         nx65922, nx65924, nx65926, nx65928, nx65930, nx65932, nx65934, nx65936, 
         nx65938, nx65940, nx65942, nx65944, nx65946, nx65948, nx65950, nx65952, 
         nx65954, nx65956, nx65958, nx65960, nx65962, nx65964, nx65966, nx65968, 
         nx65970, nx65972, nx65974, nx65976, nx65978, nx65982, nx65984, nx65986, 
         nx65988, nx65990, nx65992, nx65994, nx65996, nx65998, nx66000, nx66002, 
         nx66004, nx66006, nx66008, nx66010, nx66012, nx66014, nx66016, nx66018, 
         nx66020, nx66022, nx66024, nx66026, nx66028, nx66030, nx66032, nx66034, 
         nx66036, nx66038, nx66040, nx66042, nx66044, nx66046, nx66048, nx66050, 
         nx66052, nx66054, nx66056, nx66058, nx66060, nx66062, nx66064, nx66066, 
         nx66068, nx66070, nx66072, nx66074, nx66076, nx66078, nx66080, nx66082, 
         nx66084, nx66086, nx66088, nx66090, nx66092, nx66094, nx66096, nx66098, 
         nx66100, nx66102, nx66104, nx66106, nx66108, nx66110, nx66112, nx66114, 
         nx66116, nx66118, nx66120, nx66122, nx66124, nx66126, nx66128, nx66130, 
         nx66132, nx66134, nx66136, nx66138, nx66140, nx66142, nx66144, nx66146, 
         nx66148, nx66150, nx66152, nx66154, nx66156, nx66158, nx66160, nx66162, 
         nx66164, nx66166, nx66168, nx66170, nx66172, nx66174, nx66176, nx66178, 
         nx66180, nx66182, nx66184, nx66186, nx66188, nx66190, nx66192, nx66194, 
         nx66196, nx66198, nx66200, nx66202, nx66204, nx66206, nx66208, nx66210, 
         nx66212, nx66214, nx66216, nx66218, nx66220, nx66222, nx66224, nx66226, 
         nx66228, nx66230, nx66232, nx66234, nx66236, nx66238, nx66240, nx66242, 
         nx66244, nx66246, nx66248, nx66250, nx66252, nx66254, nx66256, nx66258, 
         nx66260, nx66262, nx66264, nx66266, nx66268, nx66270, nx66272, nx66274, 
         nx66276, nx66278, nx66280, nx66282, nx66284, nx66286;
    wire [2047:0] \$dummy ;




    or04 ix4797 (.Y (dataout[0]), .A0 (nx4792), .A1 (nx3612), .A2 (nx2436), .A3 (
         nx1256)) ;
    nand04 ix4793 (.Y (nx4792), .A0 (nx54112), .A1 (nx54273), .A2 (nx54364), .A3 (
           nx54455)) ;
    oai21 ix54113 (.Y (nx54112), .A0 (nx4782), .A1 (nx4640), .B0 (nx65096)) ;
    nand04 ix4783 (.Y (nx4782), .A0 (nx54115), .A1 (nx54142), .A2 (nx54163), .A3 (
           nx54183)) ;
    aoi22 ix54116 (.Y (nx54115), .A0 (ram_240__0), .A1 (nx64488), .B0 (
          ram_241__0), .B1 (nx65330)) ;
    dffr reg_ram_240__0 (.Q (ram_240__0), .QB (\$dummy [0]), .D (nx36180), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36181 (.Y (nx36180), .A0 (ram_240__0), .A1 (nx65982), .S0 (
             nx64414)) ;
    nand04 ix4499 (.Y (nx4498), .A0 (address[6]), .A1 (address[7]), .A2 (
           address[4]), .A3 (nx65440)) ;
    nor02_2x ix54125 (.Y (nx54124), .A0 (address[2]), .A1 (address[3])) ;
    nor02_2x ix54127 (.Y (nx54126), .A0 (address[0]), .A1 (nx65444)) ;
    nor04 ix54130 (.Y (nx54129), .A0 (address[2]), .A1 (address[3]), .A2 (
          address[0]), .A3 (nx65444)) ;
    dffr reg_ram_241__0 (.Q (ram_241__0), .QB (\$dummy [1]), .D (nx36170), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36171 (.Y (nx36170), .A0 (ram_241__0), .A1 (nx65982), .S0 (
             nx64410)) ;
    nand02 ix319 (.Y (nx318), .A0 (nx54135), .A1 (nx54124)) ;
    aoi22 ix54143 (.Y (nx54142), .A0 (ram_243__0), .A1 (nx65332), .B0 (
          ram_242__0), .B1 (nx65334)) ;
    dffr reg_ram_243__0 (.Q (ram_243__0), .QB (\$dummy [2]), .D (nx36150), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36151 (.Y (nx36150), .A0 (ram_243__0), .A1 (nx65982), .S0 (
             nx64402)) ;
    nand03 ix281 (.Y (nx280), .A0 (address[0]), .A1 (nx65444), .A2 (nx54124)) ;
    dffr reg_ram_242__0 (.Q (ram_242__0), .QB (\$dummy [3]), .D (nx36160), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36161 (.Y (nx36160), .A0 (ram_242__0), .A1 (nx65982), .S0 (
             nx64406)) ;
    nand02 ix299 (.Y (nx298), .A0 (nx54156), .A1 (nx54124)) ;
    aoi22 ix54164 (.Y (nx54163), .A0 (ram_244__0), .A1 (nx65336), .B0 (
          ram_245__0), .B1 (nx65338)) ;
    dffr reg_ram_244__0 (.Q (ram_244__0), .QB (\$dummy [4]), .D (nx36140), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36141 (.Y (nx36140), .A0 (ram_244__0), .A1 (nx65982), .S0 (
             nx64398)) ;
    nand02 ix257 (.Y (nx256), .A0 (nx54169), .A1 (nx54126)) ;
    dffr reg_ram_245__0 (.Q (ram_245__0), .QB (\$dummy [5]), .D (nx36130), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36131 (.Y (nx36130), .A0 (ram_245__0), .A1 (nx65982), .S0 (
             nx64394)) ;
    nand02 ix239 (.Y (nx238), .A0 (nx54169), .A1 (nx54135)) ;
    aoi22 ix54184 (.Y (nx54183), .A0 (ram_247__0), .A1 (nx65340), .B0 (
          ram_246__0), .B1 (nx65342)) ;
    dffr reg_ram_247__0 (.Q (ram_247__0), .QB (\$dummy [6]), .D (nx36110), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36111 (.Y (nx36110), .A0 (ram_247__0), .A1 (nx65982), .S0 (
             nx64386)) ;
    nand03 ix201 (.Y (nx200), .A0 (nx54169), .A1 (address[0]), .A2 (nx65444)) ;
    dffr reg_ram_246__0 (.Q (ram_246__0), .QB (\$dummy [7]), .D (nx36120), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36121 (.Y (nx36120), .A0 (ram_246__0), .A1 (nx65984), .S0 (
             nx64390)) ;
    nand02 ix219 (.Y (nx218), .A0 (nx54169), .A1 (nx54156)) ;
    nand04 ix4641 (.Y (nx4640), .A0 (nx54200), .A1 (nx54220), .A2 (nx54236), .A3 (
           nx54253)) ;
    aoi22 ix54201 (.Y (nx54200), .A0 (ram_248__0), .A1 (nx65344), .B0 (
          ram_249__0), .B1 (nx65346)) ;
    dffr reg_ram_248__0 (.Q (ram_248__0), .QB (\$dummy [8]), .D (nx36100), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36101 (.Y (nx36100), .A0 (ram_248__0), .A1 (nx65984), .S0 (
             nx64382)) ;
    nand02 ix173 (.Y (nx172), .A0 (nx54206), .A1 (nx54126)) ;
    dffr reg_ram_249__0 (.Q (ram_249__0), .QB (\$dummy [9]), .D (nx36090), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36091 (.Y (nx36090), .A0 (ram_249__0), .A1 (nx65984), .S0 (
             nx64378)) ;
    nand02 ix155 (.Y (nx154), .A0 (nx54206), .A1 (nx54135)) ;
    aoi22 ix54221 (.Y (nx54220), .A0 (ram_251__0), .A1 (nx65348), .B0 (
          ram_250__0), .B1 (nx65350)) ;
    dffr reg_ram_251__0 (.Q (ram_251__0), .QB (\$dummy [10]), .D (nx36070), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36071 (.Y (nx36070), .A0 (ram_251__0), .A1 (nx65984), .S0 (
             nx64370)) ;
    nand03 ix117 (.Y (nx116), .A0 (nx54206), .A1 (address[0]), .A2 (nx65444)) ;
    dffr reg_ram_250__0 (.Q (ram_250__0), .QB (\$dummy [11]), .D (nx36080), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36081 (.Y (nx36080), .A0 (ram_250__0), .A1 (nx65984), .S0 (
             nx64374)) ;
    nand02 ix135 (.Y (nx134), .A0 (nx54206), .A1 (nx54156)) ;
    aoi22 ix54237 (.Y (nx54236), .A0 (ram_252__0), .A1 (nx65352), .B0 (
          ram_253__0), .B1 (nx65354)) ;
    dffr reg_ram_252__0 (.Q (ram_252__0), .QB (\$dummy [12]), .D (nx36060), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36061 (.Y (nx36060), .A0 (ram_252__0), .A1 (nx65984), .S0 (
             nx64366)) ;
    nand03 ix91 (.Y (nx90), .A0 (address[2]), .A1 (address[3]), .A2 (nx54126)) ;
    dffr reg_ram_253__0 (.Q (ram_253__0), .QB (\$dummy [13]), .D (nx36050), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36051 (.Y (nx36050), .A0 (ram_253__0), .A1 (nx65984), .S0 (
             nx64362)) ;
    nand03 ix71 (.Y (nx70), .A0 (address[2]), .A1 (address[3]), .A2 (nx54135)) ;
    aoi22 ix54254 (.Y (nx54253), .A0 (ram_255__0), .A1 (nx65356), .B0 (
          ram_254__0), .B1 (nx65358)) ;
    dffr reg_ram_255__0 (.Q (ram_255__0), .QB (\$dummy [14]), .D (nx36030), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36031 (.Y (nx36030), .A0 (ram_255__0), .A1 (nx65986), .S0 (
             nx64354)) ;
    nand04 ix25 (.Y (nx24), .A0 (address[2]), .A1 (address[3]), .A2 (address[0])
           , .A3 (nx65444)) ;
    dffr reg_ram_254__0 (.Q (ram_254__0), .QB (\$dummy [15]), .D (nx36040), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36041 (.Y (nx36040), .A0 (ram_254__0), .A1 (nx65986), .S0 (
             nx64358)) ;
    nand03 ix47 (.Y (nx46), .A0 (address[2]), .A1 (address[3]), .A2 (nx54156)) ;
    oai21 ix54274 (.Y (nx54273), .A0 (nx4490), .A1 (nx4348), .B0 (nx65100)) ;
    nand04 ix4491 (.Y (nx4490), .A0 (nx54276), .A1 (nx54291), .A2 (nx54301), .A3 (
           nx54311)) ;
    aoi22 ix54277 (.Y (nx54276), .A0 (ram_224__0), .A1 (nx64488), .B0 (
          ram_225__0), .B1 (nx65330)) ;
    dffr reg_ram_224__0 (.Q (ram_224__0), .QB (\$dummy [16]), .D (nx36020), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36021 (.Y (nx36020), .A0 (ram_224__0), .A1 (nx65986), .S0 (
             nx64344)) ;
    nand03 ix4207 (.Y (nx4206), .A0 (address[6]), .A1 (address[7]), .A2 (nx54282
           )) ;
    dffr reg_ram_225__0 (.Q (ram_225__0), .QB (\$dummy [17]), .D (nx36010), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36011 (.Y (nx36010), .A0 (ram_225__0), .A1 (nx65986), .S0 (
             nx64340)) ;
    aoi22 ix54292 (.Y (nx54291), .A0 (ram_227__0), .A1 (nx65332), .B0 (
          ram_226__0), .B1 (nx65334)) ;
    dffr reg_ram_227__0 (.Q (ram_227__0), .QB (\$dummy [18]), .D (nx35990), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35991 (.Y (nx35990), .A0 (ram_227__0), .A1 (nx65986), .S0 (
             nx64332)) ;
    dffr reg_ram_226__0 (.Q (ram_226__0), .QB (\$dummy [19]), .D (nx36000), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36001 (.Y (nx36000), .A0 (ram_226__0), .A1 (nx65986), .S0 (
             nx64336)) ;
    aoi22 ix54302 (.Y (nx54301), .A0 (ram_228__0), .A1 (nx65336), .B0 (
          ram_229__0), .B1 (nx65338)) ;
    dffr reg_ram_228__0 (.Q (ram_228__0), .QB (\$dummy [20]), .D (nx35980), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35981 (.Y (nx35980), .A0 (ram_228__0), .A1 (nx65986), .S0 (
             nx64328)) ;
    dffr reg_ram_229__0 (.Q (ram_229__0), .QB (\$dummy [21]), .D (nx35970), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35971 (.Y (nx35970), .A0 (ram_229__0), .A1 (nx65988), .S0 (
             nx64324)) ;
    aoi22 ix54312 (.Y (nx54311), .A0 (ram_231__0), .A1 (nx65340), .B0 (
          ram_230__0), .B1 (nx65342)) ;
    dffr reg_ram_231__0 (.Q (ram_231__0), .QB (\$dummy [22]), .D (nx35950), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35951 (.Y (nx35950), .A0 (ram_231__0), .A1 (nx65988), .S0 (
             nx64316)) ;
    dffr reg_ram_230__0 (.Q (ram_230__0), .QB (\$dummy [23]), .D (nx35960), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35961 (.Y (nx35960), .A0 (ram_230__0), .A1 (nx65988), .S0 (
             nx64320)) ;
    nand04 ix4349 (.Y (nx4348), .A0 (nx54322), .A1 (nx54332), .A2 (nx54342), .A3 (
           nx54352)) ;
    aoi22 ix54323 (.Y (nx54322), .A0 (ram_232__0), .A1 (nx65344), .B0 (
          ram_233__0), .B1 (nx65346)) ;
    dffr reg_ram_232__0 (.Q (ram_232__0), .QB (\$dummy [24]), .D (nx35940), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35941 (.Y (nx35940), .A0 (ram_232__0), .A1 (nx65988), .S0 (
             nx64312)) ;
    dffr reg_ram_233__0 (.Q (ram_233__0), .QB (\$dummy [25]), .D (nx35930), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35931 (.Y (nx35930), .A0 (ram_233__0), .A1 (nx65988), .S0 (
             nx64308)) ;
    aoi22 ix54333 (.Y (nx54332), .A0 (ram_235__0), .A1 (nx65348), .B0 (
          ram_234__0), .B1 (nx65350)) ;
    dffr reg_ram_235__0 (.Q (ram_235__0), .QB (\$dummy [26]), .D (nx35910), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35911 (.Y (nx35910), .A0 (ram_235__0), .A1 (nx65988), .S0 (
             nx64300)) ;
    dffr reg_ram_234__0 (.Q (ram_234__0), .QB (\$dummy [27]), .D (nx35920), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35921 (.Y (nx35920), .A0 (ram_234__0), .A1 (nx65988), .S0 (
             nx64304)) ;
    aoi22 ix54343 (.Y (nx54342), .A0 (ram_236__0), .A1 (nx65352), .B0 (
          ram_237__0), .B1 (nx65354)) ;
    dffr reg_ram_236__0 (.Q (ram_236__0), .QB (\$dummy [28]), .D (nx35900), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35901 (.Y (nx35900), .A0 (ram_236__0), .A1 (nx65990), .S0 (
             nx64296)) ;
    dffr reg_ram_237__0 (.Q (ram_237__0), .QB (\$dummy [29]), .D (nx35890), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35891 (.Y (nx35890), .A0 (ram_237__0), .A1 (nx65990), .S0 (
             nx64292)) ;
    aoi22 ix54353 (.Y (nx54352), .A0 (ram_239__0), .A1 (nx65356), .B0 (
          ram_238__0), .B1 (nx65358)) ;
    dffr reg_ram_239__0 (.Q (ram_239__0), .QB (\$dummy [30]), .D (nx35870), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35871 (.Y (nx35870), .A0 (ram_239__0), .A1 (nx65990), .S0 (
             nx64284)) ;
    dffr reg_ram_238__0 (.Q (ram_238__0), .QB (\$dummy [31]), .D (nx35880), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35881 (.Y (nx35880), .A0 (ram_238__0), .A1 (nx65990), .S0 (
             nx64288)) ;
    oai21 ix54365 (.Y (nx54364), .A0 (nx4196), .A1 (nx4054), .B0 (nx65104)) ;
    nand04 ix4197 (.Y (nx4196), .A0 (nx54367), .A1 (nx54382), .A2 (nx54392), .A3 (
           nx54402)) ;
    aoi22 ix54368 (.Y (nx54367), .A0 (ram_208__0), .A1 (nx64488), .B0 (
          ram_209__0), .B1 (nx65330)) ;
    dffr reg_ram_208__0 (.Q (ram_208__0), .QB (\$dummy [32]), .D (nx35860), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35861 (.Y (nx35860), .A0 (ram_208__0), .A1 (nx65990), .S0 (
             nx64274)) ;
    nand03 ix3913 (.Y (nx3912), .A0 (address[6]), .A1 (address[7]), .A2 (nx54373
           )) ;
    dffr reg_ram_209__0 (.Q (ram_209__0), .QB (\$dummy [33]), .D (nx35850), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35851 (.Y (nx35850), .A0 (ram_209__0), .A1 (nx65990), .S0 (
             nx64270)) ;
    aoi22 ix54383 (.Y (nx54382), .A0 (ram_211__0), .A1 (nx65332), .B0 (
          ram_210__0), .B1 (nx65334)) ;
    dffr reg_ram_211__0 (.Q (ram_211__0), .QB (\$dummy [34]), .D (nx35830), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35831 (.Y (nx35830), .A0 (ram_211__0), .A1 (nx65990), .S0 (
             nx64262)) ;
    dffr reg_ram_210__0 (.Q (ram_210__0), .QB (\$dummy [35]), .D (nx35840), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35841 (.Y (nx35840), .A0 (ram_210__0), .A1 (nx65992), .S0 (
             nx64266)) ;
    aoi22 ix54393 (.Y (nx54392), .A0 (ram_212__0), .A1 (nx65336), .B0 (
          ram_213__0), .B1 (nx65338)) ;
    dffr reg_ram_212__0 (.Q (ram_212__0), .QB (\$dummy [36]), .D (nx35820), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35821 (.Y (nx35820), .A0 (ram_212__0), .A1 (nx65992), .S0 (
             nx64258)) ;
    dffr reg_ram_213__0 (.Q (ram_213__0), .QB (\$dummy [37]), .D (nx35810), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35811 (.Y (nx35810), .A0 (ram_213__0), .A1 (nx65992), .S0 (
             nx64254)) ;
    aoi22 ix54403 (.Y (nx54402), .A0 (ram_215__0), .A1 (nx65340), .B0 (
          ram_214__0), .B1 (nx65342)) ;
    dffr reg_ram_215__0 (.Q (ram_215__0), .QB (\$dummy [38]), .D (nx35790), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35791 (.Y (nx35790), .A0 (ram_215__0), .A1 (nx65992), .S0 (
             nx64246)) ;
    dffr reg_ram_214__0 (.Q (ram_214__0), .QB (\$dummy [39]), .D (nx35800), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35801 (.Y (nx35800), .A0 (ram_214__0), .A1 (nx65992), .S0 (
             nx64250)) ;
    nand04 ix4055 (.Y (nx4054), .A0 (nx54413), .A1 (nx54423), .A2 (nx54433), .A3 (
           nx54443)) ;
    aoi22 ix54414 (.Y (nx54413), .A0 (ram_216__0), .A1 (nx65344), .B0 (
          ram_217__0), .B1 (nx65346)) ;
    dffr reg_ram_216__0 (.Q (ram_216__0), .QB (\$dummy [40]), .D (nx35780), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35781 (.Y (nx35780), .A0 (ram_216__0), .A1 (nx65992), .S0 (
             nx64242)) ;
    dffr reg_ram_217__0 (.Q (ram_217__0), .QB (\$dummy [41]), .D (nx35770), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35771 (.Y (nx35770), .A0 (ram_217__0), .A1 (nx65992), .S0 (
             nx64238)) ;
    aoi22 ix54424 (.Y (nx54423), .A0 (ram_219__0), .A1 (nx65348), .B0 (
          ram_218__0), .B1 (nx65350)) ;
    dffr reg_ram_219__0 (.Q (ram_219__0), .QB (\$dummy [42]), .D (nx35750), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35751 (.Y (nx35750), .A0 (ram_219__0), .A1 (nx65994), .S0 (
             nx64230)) ;
    dffr reg_ram_218__0 (.Q (ram_218__0), .QB (\$dummy [43]), .D (nx35760), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35761 (.Y (nx35760), .A0 (ram_218__0), .A1 (nx65994), .S0 (
             nx64234)) ;
    aoi22 ix54434 (.Y (nx54433), .A0 (ram_220__0), .A1 (nx65352), .B0 (
          ram_221__0), .B1 (nx65354)) ;
    dffr reg_ram_220__0 (.Q (ram_220__0), .QB (\$dummy [44]), .D (nx35740), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35741 (.Y (nx35740), .A0 (ram_220__0), .A1 (nx65994), .S0 (
             nx64226)) ;
    dffr reg_ram_221__0 (.Q (ram_221__0), .QB (\$dummy [45]), .D (nx35730), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35731 (.Y (nx35730), .A0 (ram_221__0), .A1 (nx65994), .S0 (
             nx64222)) ;
    aoi22 ix54444 (.Y (nx54443), .A0 (ram_223__0), .A1 (nx65356), .B0 (
          ram_222__0), .B1 (nx65358)) ;
    dffr reg_ram_223__0 (.Q (ram_223__0), .QB (\$dummy [46]), .D (nx35710), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35711 (.Y (nx35710), .A0 (ram_223__0), .A1 (nx65994), .S0 (
             nx64214)) ;
    dffr reg_ram_222__0 (.Q (ram_222__0), .QB (\$dummy [47]), .D (nx35720), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35721 (.Y (nx35720), .A0 (ram_222__0), .A1 (nx65994), .S0 (
             nx64218)) ;
    oai21 ix54456 (.Y (nx54455), .A0 (nx3904), .A1 (nx3762), .B0 (nx65108)) ;
    nand04 ix3905 (.Y (nx3904), .A0 (nx54458), .A1 (nx54471), .A2 (nx54481), .A3 (
           nx54491)) ;
    aoi22 ix54459 (.Y (nx54458), .A0 (ram_192__0), .A1 (nx64488), .B0 (
          ram_193__0), .B1 (nx65330)) ;
    dffr reg_ram_192__0 (.Q (ram_192__0), .QB (\$dummy [48]), .D (nx35700), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35701 (.Y (nx35700), .A0 (ram_192__0), .A1 (nx65994), .S0 (
             nx64204)) ;
    nand03 ix3621 (.Y (nx3620), .A0 (address[6]), .A1 (address[7]), .A2 (nx54464
           )) ;
    nor02_2x ix54465 (.Y (nx54464), .A0 (address[4]), .A1 (nx65440)) ;
    dffr reg_ram_193__0 (.Q (ram_193__0), .QB (\$dummy [49]), .D (nx35690), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35691 (.Y (nx35690), .A0 (ram_193__0), .A1 (nx65996), .S0 (
             nx64200)) ;
    aoi22 ix54472 (.Y (nx54471), .A0 (ram_195__0), .A1 (nx65332), .B0 (
          ram_194__0), .B1 (nx65334)) ;
    dffr reg_ram_195__0 (.Q (ram_195__0), .QB (\$dummy [50]), .D (nx35670), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35671 (.Y (nx35670), .A0 (ram_195__0), .A1 (nx65996), .S0 (
             nx64192)) ;
    dffr reg_ram_194__0 (.Q (ram_194__0), .QB (\$dummy [51]), .D (nx35680), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35681 (.Y (nx35680), .A0 (ram_194__0), .A1 (nx65996), .S0 (
             nx64196)) ;
    aoi22 ix54482 (.Y (nx54481), .A0 (ram_196__0), .A1 (nx65336), .B0 (
          ram_197__0), .B1 (nx65338)) ;
    dffr reg_ram_196__0 (.Q (ram_196__0), .QB (\$dummy [52]), .D (nx35660), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35661 (.Y (nx35660), .A0 (ram_196__0), .A1 (nx65996), .S0 (
             nx64188)) ;
    dffr reg_ram_197__0 (.Q (ram_197__0), .QB (\$dummy [53]), .D (nx35650), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35651 (.Y (nx35650), .A0 (ram_197__0), .A1 (nx65996), .S0 (
             nx64184)) ;
    aoi22 ix54492 (.Y (nx54491), .A0 (ram_199__0), .A1 (nx65340), .B0 (
          ram_198__0), .B1 (nx65342)) ;
    dffr reg_ram_199__0 (.Q (ram_199__0), .QB (\$dummy [54]), .D (nx35630), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35631 (.Y (nx35630), .A0 (ram_199__0), .A1 (nx65996), .S0 (
             nx64176)) ;
    dffr reg_ram_198__0 (.Q (ram_198__0), .QB (\$dummy [55]), .D (nx35640), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35641 (.Y (nx35640), .A0 (ram_198__0), .A1 (nx65996), .S0 (
             nx64180)) ;
    nand04 ix3763 (.Y (nx3762), .A0 (nx54502), .A1 (nx54512), .A2 (nx54522), .A3 (
           nx54532)) ;
    aoi22 ix54503 (.Y (nx54502), .A0 (ram_200__0), .A1 (nx65344), .B0 (
          ram_201__0), .B1 (nx65346)) ;
    dffr reg_ram_200__0 (.Q (ram_200__0), .QB (\$dummy [56]), .D (nx35620), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35621 (.Y (nx35620), .A0 (ram_200__0), .A1 (nx65998), .S0 (
             nx64172)) ;
    dffr reg_ram_201__0 (.Q (ram_201__0), .QB (\$dummy [57]), .D (nx35610), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35611 (.Y (nx35610), .A0 (ram_201__0), .A1 (nx65998), .S0 (
             nx64168)) ;
    aoi22 ix54513 (.Y (nx54512), .A0 (ram_203__0), .A1 (nx65348), .B0 (
          ram_202__0), .B1 (nx65350)) ;
    dffr reg_ram_203__0 (.Q (ram_203__0), .QB (\$dummy [58]), .D (nx35590), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35591 (.Y (nx35590), .A0 (ram_203__0), .A1 (nx65998), .S0 (
             nx64160)) ;
    dffr reg_ram_202__0 (.Q (ram_202__0), .QB (\$dummy [59]), .D (nx35600), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35601 (.Y (nx35600), .A0 (ram_202__0), .A1 (nx65998), .S0 (
             nx64164)) ;
    aoi22 ix54523 (.Y (nx54522), .A0 (ram_204__0), .A1 (nx65352), .B0 (
          ram_205__0), .B1 (nx65354)) ;
    dffr reg_ram_204__0 (.Q (ram_204__0), .QB (\$dummy [60]), .D (nx35580), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35581 (.Y (nx35580), .A0 (ram_204__0), .A1 (nx65998), .S0 (
             nx64156)) ;
    dffr reg_ram_205__0 (.Q (ram_205__0), .QB (\$dummy [61]), .D (nx35570), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35571 (.Y (nx35570), .A0 (ram_205__0), .A1 (nx65998), .S0 (
             nx64152)) ;
    aoi22 ix54533 (.Y (nx54532), .A0 (ram_207__0), .A1 (nx65356), .B0 (
          ram_206__0), .B1 (nx65358)) ;
    dffr reg_ram_207__0 (.Q (ram_207__0), .QB (\$dummy [62]), .D (nx35550), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35551 (.Y (nx35550), .A0 (ram_207__0), .A1 (nx65998), .S0 (
             nx64144)) ;
    dffr reg_ram_206__0 (.Q (ram_206__0), .QB (\$dummy [63]), .D (nx35560), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35561 (.Y (nx35560), .A0 (ram_206__0), .A1 (nx66000), .S0 (
             nx64148)) ;
    nand04 ix3613 (.Y (nx3612), .A0 (nx54545), .A1 (nx54636), .A2 (nx54723), .A3 (
           nx54812)) ;
    oai21 ix54546 (.Y (nx54545), .A0 (nx3602), .A1 (nx3460), .B0 (nx65112)) ;
    nand04 ix3603 (.Y (nx3602), .A0 (nx54548), .A1 (nx54563), .A2 (nx54573), .A3 (
           nx54583)) ;
    aoi22 ix54549 (.Y (nx54548), .A0 (ram_80__0), .A1 (nx64488), .B0 (ram_81__0)
          , .B1 (nx65330)) ;
    dffr reg_ram_80__0 (.Q (ram_80__0), .QB (\$dummy [64]), .D (nx35540), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35541 (.Y (nx35540), .A0 (ram_80__0), .A1 (nx66000), .S0 (nx64134
             )) ;
    nand02 ix3319 (.Y (nx3318), .A0 (nx54554), .A1 (nx54373)) ;
    dffr reg_ram_81__0 (.Q (ram_81__0), .QB (\$dummy [65]), .D (nx35530), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35531 (.Y (nx35530), .A0 (ram_81__0), .A1 (nx66000), .S0 (nx64130
             )) ;
    aoi22 ix54564 (.Y (nx54563), .A0 (ram_83__0), .A1 (nx65332), .B0 (ram_82__0)
          , .B1 (nx65334)) ;
    dffr reg_ram_83__0 (.Q (ram_83__0), .QB (\$dummy [66]), .D (nx35510), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35511 (.Y (nx35510), .A0 (ram_83__0), .A1 (nx66000), .S0 (nx64122
             )) ;
    dffr reg_ram_82__0 (.Q (ram_82__0), .QB (\$dummy [67]), .D (nx35520), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35521 (.Y (nx35520), .A0 (ram_82__0), .A1 (nx66000), .S0 (nx64126
             )) ;
    aoi22 ix54574 (.Y (nx54573), .A0 (ram_84__0), .A1 (nx65336), .B0 (ram_85__0)
          , .B1 (nx65338)) ;
    dffr reg_ram_84__0 (.Q (ram_84__0), .QB (\$dummy [68]), .D (nx35500), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35501 (.Y (nx35500), .A0 (ram_84__0), .A1 (nx66000), .S0 (nx64118
             )) ;
    dffr reg_ram_85__0 (.Q (ram_85__0), .QB (\$dummy [69]), .D (nx35490), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35491 (.Y (nx35490), .A0 (ram_85__0), .A1 (nx66000), .S0 (nx64114
             )) ;
    aoi22 ix54584 (.Y (nx54583), .A0 (ram_87__0), .A1 (nx65340), .B0 (ram_86__0)
          , .B1 (nx65342)) ;
    dffr reg_ram_87__0 (.Q (ram_87__0), .QB (\$dummy [70]), .D (nx35470), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35471 (.Y (nx35470), .A0 (ram_87__0), .A1 (nx66002), .S0 (nx64106
             )) ;
    dffr reg_ram_86__0 (.Q (ram_86__0), .QB (\$dummy [71]), .D (nx35480), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35481 (.Y (nx35480), .A0 (ram_86__0), .A1 (nx66002), .S0 (nx64110
             )) ;
    nand04 ix3461 (.Y (nx3460), .A0 (nx54594), .A1 (nx54604), .A2 (nx54614), .A3 (
           nx54624)) ;
    aoi22 ix54595 (.Y (nx54594), .A0 (ram_88__0), .A1 (nx65344), .B0 (ram_89__0)
          , .B1 (nx65346)) ;
    dffr reg_ram_88__0 (.Q (ram_88__0), .QB (\$dummy [72]), .D (nx35460), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35461 (.Y (nx35460), .A0 (ram_88__0), .A1 (nx66002), .S0 (nx64102
             )) ;
    dffr reg_ram_89__0 (.Q (ram_89__0), .QB (\$dummy [73]), .D (nx35450), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35451 (.Y (nx35450), .A0 (ram_89__0), .A1 (nx66002), .S0 (nx64098
             )) ;
    aoi22 ix54605 (.Y (nx54604), .A0 (ram_91__0), .A1 (nx65348), .B0 (ram_90__0)
          , .B1 (nx65350)) ;
    dffr reg_ram_91__0 (.Q (ram_91__0), .QB (\$dummy [74]), .D (nx35430), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35431 (.Y (nx35430), .A0 (ram_91__0), .A1 (nx66002), .S0 (nx64090
             )) ;
    dffr reg_ram_90__0 (.Q (ram_90__0), .QB (\$dummy [75]), .D (nx35440), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35441 (.Y (nx35440), .A0 (ram_90__0), .A1 (nx66002), .S0 (nx64094
             )) ;
    aoi22 ix54615 (.Y (nx54614), .A0 (ram_92__0), .A1 (nx65352), .B0 (ram_93__0)
          , .B1 (nx65354)) ;
    dffr reg_ram_92__0 (.Q (ram_92__0), .QB (\$dummy [76]), .D (nx35420), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35421 (.Y (nx35420), .A0 (ram_92__0), .A1 (nx66002), .S0 (nx64086
             )) ;
    dffr reg_ram_93__0 (.Q (ram_93__0), .QB (\$dummy [77]), .D (nx35410), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35411 (.Y (nx35410), .A0 (ram_93__0), .A1 (nx66004), .S0 (nx64082
             )) ;
    aoi22 ix54625 (.Y (nx54624), .A0 (ram_95__0), .A1 (nx65356), .B0 (ram_94__0)
          , .B1 (nx65358)) ;
    dffr reg_ram_95__0 (.Q (ram_95__0), .QB (\$dummy [78]), .D (nx35390), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35391 (.Y (nx35390), .A0 (ram_95__0), .A1 (nx66004), .S0 (nx64074
             )) ;
    dffr reg_ram_94__0 (.Q (ram_94__0), .QB (\$dummy [79]), .D (nx35400), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35401 (.Y (nx35400), .A0 (ram_94__0), .A1 (nx66004), .S0 (nx64078
             )) ;
    oai21 ix54637 (.Y (nx54636), .A0 (nx3310), .A1 (nx3168), .B0 (nx65116)) ;
    nand04 ix3311 (.Y (nx3310), .A0 (nx54639), .A1 (nx54650), .A2 (nx54660), .A3 (
           nx54670)) ;
    aoi22 ix54640 (.Y (nx54639), .A0 (ram_64__0), .A1 (nx64488), .B0 (ram_65__0)
          , .B1 (nx65330)) ;
    dffr reg_ram_64__0 (.Q (ram_64__0), .QB (\$dummy [80]), .D (nx35380), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35381 (.Y (nx35380), .A0 (ram_64__0), .A1 (nx66004), .S0 (nx64064
             )) ;
    nand02 ix3027 (.Y (nx3026), .A0 (nx54554), .A1 (nx54464)) ;
    dffr reg_ram_65__0 (.Q (ram_65__0), .QB (\$dummy [81]), .D (nx35370), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35371 (.Y (nx35370), .A0 (ram_65__0), .A1 (nx66004), .S0 (nx64060
             )) ;
    aoi22 ix54651 (.Y (nx54650), .A0 (ram_67__0), .A1 (nx65332), .B0 (ram_66__0)
          , .B1 (nx65334)) ;
    dffr reg_ram_67__0 (.Q (ram_67__0), .QB (\$dummy [82]), .D (nx35350), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35351 (.Y (nx35350), .A0 (ram_67__0), .A1 (nx66004), .S0 (nx64052
             )) ;
    dffr reg_ram_66__0 (.Q (ram_66__0), .QB (\$dummy [83]), .D (nx35360), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35361 (.Y (nx35360), .A0 (ram_66__0), .A1 (nx66004), .S0 (nx64056
             )) ;
    aoi22 ix54661 (.Y (nx54660), .A0 (ram_68__0), .A1 (nx65336), .B0 (ram_69__0)
          , .B1 (nx65338)) ;
    dffr reg_ram_68__0 (.Q (ram_68__0), .QB (\$dummy [84]), .D (nx35340), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35341 (.Y (nx35340), .A0 (ram_68__0), .A1 (nx66006), .S0 (nx64048
             )) ;
    dffr reg_ram_69__0 (.Q (ram_69__0), .QB (\$dummy [85]), .D (nx35330), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35331 (.Y (nx35330), .A0 (ram_69__0), .A1 (nx66006), .S0 (nx64044
             )) ;
    aoi22 ix54671 (.Y (nx54670), .A0 (ram_71__0), .A1 (nx65340), .B0 (ram_70__0)
          , .B1 (nx65342)) ;
    dffr reg_ram_71__0 (.Q (ram_71__0), .QB (\$dummy [86]), .D (nx35310), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35311 (.Y (nx35310), .A0 (ram_71__0), .A1 (nx66006), .S0 (nx64036
             )) ;
    dffr reg_ram_70__0 (.Q (ram_70__0), .QB (\$dummy [87]), .D (nx35320), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35321 (.Y (nx35320), .A0 (ram_70__0), .A1 (nx66006), .S0 (nx64040
             )) ;
    nand04 ix3169 (.Y (nx3168), .A0 (nx54681), .A1 (nx54691), .A2 (nx54701), .A3 (
           nx54711)) ;
    aoi22 ix54682 (.Y (nx54681), .A0 (ram_72__0), .A1 (nx65344), .B0 (ram_73__0)
          , .B1 (nx65346)) ;
    dffr reg_ram_72__0 (.Q (ram_72__0), .QB (\$dummy [88]), .D (nx35300), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35301 (.Y (nx35300), .A0 (ram_72__0), .A1 (nx66006), .S0 (nx64032
             )) ;
    dffr reg_ram_73__0 (.Q (ram_73__0), .QB (\$dummy [89]), .D (nx35290), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35291 (.Y (nx35290), .A0 (ram_73__0), .A1 (nx66006), .S0 (nx64028
             )) ;
    aoi22 ix54692 (.Y (nx54691), .A0 (ram_75__0), .A1 (nx65348), .B0 (ram_74__0)
          , .B1 (nx65350)) ;
    dffr reg_ram_75__0 (.Q (ram_75__0), .QB (\$dummy [90]), .D (nx35270), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35271 (.Y (nx35270), .A0 (ram_75__0), .A1 (nx66006), .S0 (nx64020
             )) ;
    dffr reg_ram_74__0 (.Q (ram_74__0), .QB (\$dummy [91]), .D (nx35280), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35281 (.Y (nx35280), .A0 (ram_74__0), .A1 (nx66008), .S0 (nx64024
             )) ;
    aoi22 ix54702 (.Y (nx54701), .A0 (ram_76__0), .A1 (nx65352), .B0 (ram_77__0)
          , .B1 (nx65354)) ;
    dffr reg_ram_76__0 (.Q (ram_76__0), .QB (\$dummy [92]), .D (nx35260), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35261 (.Y (nx35260), .A0 (ram_76__0), .A1 (nx66008), .S0 (nx64016
             )) ;
    dffr reg_ram_77__0 (.Q (ram_77__0), .QB (\$dummy [93]), .D (nx35250), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35251 (.Y (nx35250), .A0 (ram_77__0), .A1 (nx66008), .S0 (nx64012
             )) ;
    aoi22 ix54712 (.Y (nx54711), .A0 (ram_79__0), .A1 (nx65356), .B0 (ram_78__0)
          , .B1 (nx65358)) ;
    dffr reg_ram_79__0 (.Q (ram_79__0), .QB (\$dummy [94]), .D (nx35230), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35231 (.Y (nx35230), .A0 (ram_79__0), .A1 (nx66008), .S0 (nx64004
             )) ;
    dffr reg_ram_78__0 (.Q (ram_78__0), .QB (\$dummy [95]), .D (nx35240), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35241 (.Y (nx35240), .A0 (ram_78__0), .A1 (nx66008), .S0 (nx64008
             )) ;
    oai21 ix54724 (.Y (nx54723), .A0 (nx3016), .A1 (nx2874), .B0 (nx65120)) ;
    nand04 ix3017 (.Y (nx3016), .A0 (nx54726), .A1 (nx54739), .A2 (nx54749), .A3 (
           nx54759)) ;
    aoi22 ix54727 (.Y (nx54726), .A0 (ram_48__0), .A1 (nx64488), .B0 (ram_49__0)
          , .B1 (nx65330)) ;
    dffr reg_ram_48__0 (.Q (ram_48__0), .QB (\$dummy [96]), .D (nx35220), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35221 (.Y (nx35220), .A0 (ram_48__0), .A1 (nx66008), .S0 (nx63994
             )) ;
    nand03 ix2733 (.Y (nx2732), .A0 (address[4]), .A1 (nx65440), .A2 (nx54732)
           ) ;
    nor02_2x ix54733 (.Y (nx54732), .A0 (address[6]), .A1 (address[7])) ;
    dffr reg_ram_49__0 (.Q (ram_49__0), .QB (\$dummy [97]), .D (nx35210), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35211 (.Y (nx35210), .A0 (ram_49__0), .A1 (nx66008), .S0 (nx63990
             )) ;
    aoi22 ix54740 (.Y (nx54739), .A0 (ram_51__0), .A1 (nx65332), .B0 (ram_50__0)
          , .B1 (nx65334)) ;
    dffr reg_ram_51__0 (.Q (ram_51__0), .QB (\$dummy [98]), .D (nx35190), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35191 (.Y (nx35190), .A0 (ram_51__0), .A1 (nx66010), .S0 (nx63982
             )) ;
    dffr reg_ram_50__0 (.Q (ram_50__0), .QB (\$dummy [99]), .D (nx35200), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35201 (.Y (nx35200), .A0 (ram_50__0), .A1 (nx66010), .S0 (nx63986
             )) ;
    aoi22 ix54750 (.Y (nx54749), .A0 (ram_52__0), .A1 (nx65336), .B0 (ram_53__0)
          , .B1 (nx65338)) ;
    dffr reg_ram_52__0 (.Q (ram_52__0), .QB (\$dummy [100]), .D (nx35180), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35181 (.Y (nx35180), .A0 (ram_52__0), .A1 (nx66010), .S0 (nx63978
             )) ;
    dffr reg_ram_53__0 (.Q (ram_53__0), .QB (\$dummy [101]), .D (nx35170), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35171 (.Y (nx35170), .A0 (ram_53__0), .A1 (nx66010), .S0 (nx63974
             )) ;
    aoi22 ix54760 (.Y (nx54759), .A0 (ram_55__0), .A1 (nx65340), .B0 (ram_54__0)
          , .B1 (nx65342)) ;
    dffr reg_ram_55__0 (.Q (ram_55__0), .QB (\$dummy [102]), .D (nx35150), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35151 (.Y (nx35150), .A0 (ram_55__0), .A1 (nx66010), .S0 (nx63966
             )) ;
    dffr reg_ram_54__0 (.Q (ram_54__0), .QB (\$dummy [103]), .D (nx35160), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35161 (.Y (nx35160), .A0 (ram_54__0), .A1 (nx66010), .S0 (nx63970
             )) ;
    nand04 ix2875 (.Y (nx2874), .A0 (nx54770), .A1 (nx54780), .A2 (nx54790), .A3 (
           nx54800)) ;
    aoi22 ix54771 (.Y (nx54770), .A0 (ram_56__0), .A1 (nx65344), .B0 (ram_57__0)
          , .B1 (nx65346)) ;
    dffr reg_ram_56__0 (.Q (ram_56__0), .QB (\$dummy [104]), .D (nx35140), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35141 (.Y (nx35140), .A0 (ram_56__0), .A1 (nx66010), .S0 (nx63962
             )) ;
    dffr reg_ram_57__0 (.Q (ram_57__0), .QB (\$dummy [105]), .D (nx35130), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35131 (.Y (nx35130), .A0 (ram_57__0), .A1 (nx66012), .S0 (nx63958
             )) ;
    aoi22 ix54781 (.Y (nx54780), .A0 (ram_59__0), .A1 (nx65348), .B0 (ram_58__0)
          , .B1 (nx65350)) ;
    dffr reg_ram_59__0 (.Q (ram_59__0), .QB (\$dummy [106]), .D (nx35110), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35111 (.Y (nx35110), .A0 (ram_59__0), .A1 (nx66012), .S0 (nx63950
             )) ;
    dffr reg_ram_58__0 (.Q (ram_58__0), .QB (\$dummy [107]), .D (nx35120), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35121 (.Y (nx35120), .A0 (ram_58__0), .A1 (nx66012), .S0 (nx63954
             )) ;
    aoi22 ix54791 (.Y (nx54790), .A0 (ram_60__0), .A1 (nx65352), .B0 (ram_61__0)
          , .B1 (nx65354)) ;
    dffr reg_ram_60__0 (.Q (ram_60__0), .QB (\$dummy [108]), .D (nx35100), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35101 (.Y (nx35100), .A0 (ram_60__0), .A1 (nx66012), .S0 (nx63946
             )) ;
    dffr reg_ram_61__0 (.Q (ram_61__0), .QB (\$dummy [109]), .D (nx35090), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35091 (.Y (nx35090), .A0 (ram_61__0), .A1 (nx66012), .S0 (nx63942
             )) ;
    aoi22 ix54801 (.Y (nx54800), .A0 (ram_63__0), .A1 (nx65356), .B0 (ram_62__0)
          , .B1 (nx65358)) ;
    dffr reg_ram_63__0 (.Q (ram_63__0), .QB (\$dummy [110]), .D (nx35070), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35071 (.Y (nx35070), .A0 (ram_63__0), .A1 (nx66012), .S0 (nx63934
             )) ;
    dffr reg_ram_62__0 (.Q (ram_62__0), .QB (\$dummy [111]), .D (nx35080), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35081 (.Y (nx35080), .A0 (ram_62__0), .A1 (nx66012), .S0 (nx63938
             )) ;
    oai21 ix54813 (.Y (nx54812), .A0 (nx2724), .A1 (nx2582), .B0 (nx65124)) ;
    nand04 ix2725 (.Y (nx2724), .A0 (nx54815), .A1 (nx54826), .A2 (nx54836), .A3 (
           nx54846)) ;
    aoi22 ix54816 (.Y (nx54815), .A0 (ram_32__0), .A1 (nx64490), .B0 (ram_33__0)
          , .B1 (nx64528)) ;
    dffr reg_ram_32__0 (.Q (ram_32__0), .QB (\$dummy [112]), .D (nx35060), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35061 (.Y (nx35060), .A0 (ram_32__0), .A1 (nx66014), .S0 (nx63924
             )) ;
    nand02 ix2441 (.Y (nx2440), .A0 (nx54282), .A1 (nx54732)) ;
    dffr reg_ram_33__0 (.Q (ram_33__0), .QB (\$dummy [113]), .D (nx35050), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35051 (.Y (nx35050), .A0 (ram_33__0), .A1 (nx66014), .S0 (nx63920
             )) ;
    aoi22 ix54827 (.Y (nx54826), .A0 (ram_35__0), .A1 (nx64566), .B0 (ram_34__0)
          , .B1 (nx64604)) ;
    dffr reg_ram_35__0 (.Q (ram_35__0), .QB (\$dummy [114]), .D (nx35030), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35031 (.Y (nx35030), .A0 (ram_35__0), .A1 (nx66014), .S0 (nx63912
             )) ;
    dffr reg_ram_34__0 (.Q (ram_34__0), .QB (\$dummy [115]), .D (nx35040), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35041 (.Y (nx35040), .A0 (ram_34__0), .A1 (nx66014), .S0 (nx63916
             )) ;
    aoi22 ix54837 (.Y (nx54836), .A0 (ram_36__0), .A1 (nx64642), .B0 (ram_37__0)
          , .B1 (nx64680)) ;
    dffr reg_ram_36__0 (.Q (ram_36__0), .QB (\$dummy [116]), .D (nx35020), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35021 (.Y (nx35020), .A0 (ram_36__0), .A1 (nx66014), .S0 (nx63908
             )) ;
    dffr reg_ram_37__0 (.Q (ram_37__0), .QB (\$dummy [117]), .D (nx35010), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35011 (.Y (nx35010), .A0 (ram_37__0), .A1 (nx66014), .S0 (nx63904
             )) ;
    aoi22 ix54847 (.Y (nx54846), .A0 (ram_39__0), .A1 (nx64718), .B0 (ram_38__0)
          , .B1 (nx64756)) ;
    dffr reg_ram_39__0 (.Q (ram_39__0), .QB (\$dummy [118]), .D (nx34990), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34991 (.Y (nx34990), .A0 (ram_39__0), .A1 (nx66014), .S0 (nx63896
             )) ;
    dffr reg_ram_38__0 (.Q (ram_38__0), .QB (\$dummy [119]), .D (nx35000), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix35001 (.Y (nx35000), .A0 (ram_38__0), .A1 (nx66016), .S0 (nx63900
             )) ;
    nand04 ix2583 (.Y (nx2582), .A0 (nx54857), .A1 (nx54867), .A2 (nx54877), .A3 (
           nx54887)) ;
    aoi22 ix54858 (.Y (nx54857), .A0 (ram_40__0), .A1 (nx64794), .B0 (ram_41__0)
          , .B1 (nx64832)) ;
    dffr reg_ram_40__0 (.Q (ram_40__0), .QB (\$dummy [120]), .D (nx34980), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34981 (.Y (nx34980), .A0 (ram_40__0), .A1 (nx66016), .S0 (nx63892
             )) ;
    dffr reg_ram_41__0 (.Q (ram_41__0), .QB (\$dummy [121]), .D (nx34970), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34971 (.Y (nx34970), .A0 (ram_41__0), .A1 (nx66016), .S0 (nx63888
             )) ;
    aoi22 ix54868 (.Y (nx54867), .A0 (ram_43__0), .A1 (nx64870), .B0 (ram_42__0)
          , .B1 (nx64908)) ;
    dffr reg_ram_43__0 (.Q (ram_43__0), .QB (\$dummy [122]), .D (nx34950), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34951 (.Y (nx34950), .A0 (ram_43__0), .A1 (nx66016), .S0 (nx63880
             )) ;
    dffr reg_ram_42__0 (.Q (ram_42__0), .QB (\$dummy [123]), .D (nx34960), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34961 (.Y (nx34960), .A0 (ram_42__0), .A1 (nx66016), .S0 (nx63884
             )) ;
    aoi22 ix54878 (.Y (nx54877), .A0 (ram_44__0), .A1 (nx64946), .B0 (ram_45__0)
          , .B1 (nx64984)) ;
    dffr reg_ram_44__0 (.Q (ram_44__0), .QB (\$dummy [124]), .D (nx34940), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34941 (.Y (nx34940), .A0 (ram_44__0), .A1 (nx66016), .S0 (nx63876
             )) ;
    dffr reg_ram_45__0 (.Q (ram_45__0), .QB (\$dummy [125]), .D (nx34930), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34931 (.Y (nx34930), .A0 (ram_45__0), .A1 (nx66016), .S0 (nx63872
             )) ;
    aoi22 ix54888 (.Y (nx54887), .A0 (ram_47__0), .A1 (nx65022), .B0 (ram_46__0)
          , .B1 (nx65060)) ;
    dffr reg_ram_47__0 (.Q (ram_47__0), .QB (\$dummy [126]), .D (nx34910), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34911 (.Y (nx34910), .A0 (ram_47__0), .A1 (nx66018), .S0 (nx63864
             )) ;
    dffr reg_ram_46__0 (.Q (ram_46__0), .QB (\$dummy [127]), .D (nx34920), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34921 (.Y (nx34920), .A0 (ram_46__0), .A1 (nx66018), .S0 (nx63868
             )) ;
    nand04 ix2437 (.Y (nx2436), .A0 (nx54900), .A1 (nx54987), .A2 (nx55089), .A3 (
           nx55176)) ;
    oai21 ix54901 (.Y (nx54900), .A0 (nx2426), .A1 (nx2284), .B0 (nx65128)) ;
    nand04 ix2427 (.Y (nx2426), .A0 (nx54903), .A1 (nx54914), .A2 (nx54924), .A3 (
           nx54934)) ;
    aoi22 ix54904 (.Y (nx54903), .A0 (ram_16__0), .A1 (nx64490), .B0 (ram_17__0)
          , .B1 (nx64528)) ;
    dffr reg_ram_16__0 (.Q (ram_16__0), .QB (\$dummy [128]), .D (nx34900), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34901 (.Y (nx34900), .A0 (ram_16__0), .A1 (nx66018), .S0 (nx63854
             )) ;
    nand02 ix2143 (.Y (nx2142), .A0 (nx54373), .A1 (nx54732)) ;
    dffr reg_ram_17__0 (.Q (ram_17__0), .QB (\$dummy [129]), .D (nx34890), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34891 (.Y (nx34890), .A0 (ram_17__0), .A1 (nx66018), .S0 (nx63850
             )) ;
    aoi22 ix54915 (.Y (nx54914), .A0 (ram_19__0), .A1 (nx64566), .B0 (ram_18__0)
          , .B1 (nx64604)) ;
    dffr reg_ram_19__0 (.Q (ram_19__0), .QB (\$dummy [130]), .D (nx34870), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34871 (.Y (nx34870), .A0 (ram_19__0), .A1 (nx66018), .S0 (nx63842
             )) ;
    dffr reg_ram_18__0 (.Q (ram_18__0), .QB (\$dummy [131]), .D (nx34880), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34881 (.Y (nx34880), .A0 (ram_18__0), .A1 (nx66018), .S0 (nx63846
             )) ;
    aoi22 ix54925 (.Y (nx54924), .A0 (ram_20__0), .A1 (nx64642), .B0 (ram_21__0)
          , .B1 (nx64680)) ;
    dffr reg_ram_20__0 (.Q (ram_20__0), .QB (\$dummy [132]), .D (nx34860), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34861 (.Y (nx34860), .A0 (ram_20__0), .A1 (nx66018), .S0 (nx63838
             )) ;
    dffr reg_ram_21__0 (.Q (ram_21__0), .QB (\$dummy [133]), .D (nx34850), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34851 (.Y (nx34850), .A0 (ram_21__0), .A1 (nx66020), .S0 (nx63834
             )) ;
    aoi22 ix54935 (.Y (nx54934), .A0 (ram_23__0), .A1 (nx64718), .B0 (ram_22__0)
          , .B1 (nx64756)) ;
    dffr reg_ram_23__0 (.Q (ram_23__0), .QB (\$dummy [134]), .D (nx34830), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34831 (.Y (nx34830), .A0 (ram_23__0), .A1 (nx66020), .S0 (nx63826
             )) ;
    dffr reg_ram_22__0 (.Q (ram_22__0), .QB (\$dummy [135]), .D (nx34840), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34841 (.Y (nx34840), .A0 (ram_22__0), .A1 (nx66020), .S0 (nx63830
             )) ;
    nand04 ix2285 (.Y (nx2284), .A0 (nx54945), .A1 (nx54955), .A2 (nx54965), .A3 (
           nx54975)) ;
    aoi22 ix54946 (.Y (nx54945), .A0 (ram_24__0), .A1 (nx64794), .B0 (ram_25__0)
          , .B1 (nx64832)) ;
    dffr reg_ram_24__0 (.Q (ram_24__0), .QB (\$dummy [136]), .D (nx34820), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34821 (.Y (nx34820), .A0 (ram_24__0), .A1 (nx66020), .S0 (nx63822
             )) ;
    dffr reg_ram_25__0 (.Q (ram_25__0), .QB (\$dummy [137]), .D (nx34810), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34811 (.Y (nx34810), .A0 (ram_25__0), .A1 (nx66020), .S0 (nx63818
             )) ;
    aoi22 ix54956 (.Y (nx54955), .A0 (ram_27__0), .A1 (nx64870), .B0 (ram_26__0)
          , .B1 (nx64908)) ;
    dffr reg_ram_27__0 (.Q (ram_27__0), .QB (\$dummy [138]), .D (nx34790), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34791 (.Y (nx34790), .A0 (ram_27__0), .A1 (nx66020), .S0 (nx63810
             )) ;
    dffr reg_ram_26__0 (.Q (ram_26__0), .QB (\$dummy [139]), .D (nx34800), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34801 (.Y (nx34800), .A0 (ram_26__0), .A1 (nx66020), .S0 (nx63814
             )) ;
    aoi22 ix54966 (.Y (nx54965), .A0 (ram_28__0), .A1 (nx64946), .B0 (ram_29__0)
          , .B1 (nx64984)) ;
    dffr reg_ram_28__0 (.Q (ram_28__0), .QB (\$dummy [140]), .D (nx34780), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34781 (.Y (nx34780), .A0 (ram_28__0), .A1 (nx66022), .S0 (nx63806
             )) ;
    dffr reg_ram_29__0 (.Q (ram_29__0), .QB (\$dummy [141]), .D (nx34770), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34771 (.Y (nx34770), .A0 (ram_29__0), .A1 (nx66022), .S0 (nx63802
             )) ;
    aoi22 ix54976 (.Y (nx54975), .A0 (ram_31__0), .A1 (nx65022), .B0 (ram_30__0)
          , .B1 (nx65060)) ;
    dffr reg_ram_31__0 (.Q (ram_31__0), .QB (\$dummy [142]), .D (nx34750), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34751 (.Y (nx34750), .A0 (ram_31__0), .A1 (nx66022), .S0 (nx63794
             )) ;
    dffr reg_ram_30__0 (.Q (ram_30__0), .QB (\$dummy [143]), .D (nx34760), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34761 (.Y (nx34760), .A0 (ram_30__0), .A1 (nx66022), .S0 (nx63798
             )) ;
    oai21 ix54988 (.Y (nx54987), .A0 (nx2134), .A1 (nx1992), .B0 (nx65142)) ;
    nand04 ix2135 (.Y (nx2134), .A0 (nx54990), .A1 (nx55004), .A2 (nx55016), .A3 (
           nx55028)) ;
    aoi22 ix54991 (.Y (nx54990), .A0 (ram_0__0), .A1 (nx64490), .B0 (ram_1__0), 
          .B1 (nx64528)) ;
    dffr reg_ram_0__0 (.Q (ram_0__0), .QB (\$dummy [144]), .D (nx34740), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34741 (.Y (nx34740), .A0 (nx66022), .A1 (ram_0__0), .S0 (nx65132)
             ) ;
    nand03 ix54995 (.Y (nx54994), .A0 (nx65138), .A1 (nx65366), .A2 (nx64490)) ;
    nor04 ix54997 (.Y (nx54996), .A0 (address[6]), .A1 (address[7]), .A2 (
          address[4]), .A3 (nx65440)) ;
    dffr reg_ram_1__0 (.Q (ram_1__0), .QB (\$dummy [145]), .D (nx34730), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34731 (.Y (nx34730), .A0 (nx66022), .A1 (ram_1__0), .S0 (nx65146)
             ) ;
    nand03 ix55002 (.Y (nx55001), .A0 (nx64528), .A1 (nx65366), .A2 (nx65138)) ;
    aoi22 ix55005 (.Y (nx55004), .A0 (ram_3__0), .A1 (nx64566), .B0 (ram_2__0), 
          .B1 (nx64604)) ;
    dffr reg_ram_3__0 (.Q (ram_3__0), .QB (\$dummy [146]), .D (nx34710), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34711 (.Y (nx34710), .A0 (nx66022), .A1 (ram_3__0), .S0 (nx65150)
             ) ;
    nand03 ix55009 (.Y (nx55008), .A0 (nx64566), .A1 (nx65366), .A2 (nx65138)) ;
    dffr reg_ram_2__0 (.Q (ram_2__0), .QB (\$dummy [147]), .D (nx34720), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34721 (.Y (nx34720), .A0 (nx66024), .A1 (ram_2__0), .S0 (nx65154)
             ) ;
    nand03 ix55014 (.Y (nx55013), .A0 (nx64604), .A1 (nx65366), .A2 (nx65138)) ;
    aoi22 ix55017 (.Y (nx55016), .A0 (ram_4__0), .A1 (nx64642), .B0 (ram_5__0), 
          .B1 (nx64680)) ;
    dffr reg_ram_4__0 (.Q (ram_4__0), .QB (\$dummy [148]), .D (nx34700), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34701 (.Y (nx34700), .A0 (nx66024), .A1 (ram_4__0), .S0 (nx65158)
             ) ;
    nand03 ix55021 (.Y (nx55020), .A0 (nx64642), .A1 (nx65366), .A2 (nx65138)) ;
    dffr reg_ram_5__0 (.Q (ram_5__0), .QB (\$dummy [149]), .D (nx34690), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34691 (.Y (nx34690), .A0 (nx66024), .A1 (ram_5__0), .S0 (nx65162)
             ) ;
    nand03 ix55026 (.Y (nx55025), .A0 (nx64680), .A1 (nx65366), .A2 (nx65138)) ;
    aoi22 ix55029 (.Y (nx55028), .A0 (ram_7__0), .A1 (nx64718), .B0 (ram_6__0), 
          .B1 (nx64756)) ;
    dffr reg_ram_7__0 (.Q (ram_7__0), .QB (\$dummy [150]), .D (nx34670), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34671 (.Y (nx34670), .A0 (nx66024), .A1 (ram_7__0), .S0 (nx65166)
             ) ;
    nand03 ix55033 (.Y (nx55032), .A0 (nx64718), .A1 (nx65366), .A2 (nx65138)) ;
    dffr reg_ram_6__0 (.Q (ram_6__0), .QB (\$dummy [151]), .D (nx34680), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34681 (.Y (nx34680), .A0 (nx66024), .A1 (ram_6__0), .S0 (nx65170)
             ) ;
    nand03 ix55038 (.Y (nx55037), .A0 (nx64756), .A1 (nx65368), .A2 (nx65140)) ;
    nand04 ix1993 (.Y (nx1992), .A0 (nx55041), .A1 (nx55053), .A2 (nx55065), .A3 (
           nx55077)) ;
    aoi22 ix55042 (.Y (nx55041), .A0 (ram_8__0), .A1 (nx64794), .B0 (ram_9__0), 
          .B1 (nx64832)) ;
    dffr reg_ram_8__0 (.Q (ram_8__0), .QB (\$dummy [152]), .D (nx34660), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34661 (.Y (nx34660), .A0 (nx66024), .A1 (ram_8__0), .S0 (nx65174)
             ) ;
    nand03 ix55046 (.Y (nx55045), .A0 (nx64794), .A1 (nx65368), .A2 (nx65140)) ;
    dffr reg_ram_9__0 (.Q (ram_9__0), .QB (\$dummy [153]), .D (nx34650), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34651 (.Y (nx34650), .A0 (nx66024), .A1 (ram_9__0), .S0 (nx65178)
             ) ;
    nand03 ix55051 (.Y (nx55050), .A0 (nx64832), .A1 (nx65368), .A2 (nx65140)) ;
    aoi22 ix55054 (.Y (nx55053), .A0 (ram_11__0), .A1 (nx64870), .B0 (ram_10__0)
          , .B1 (nx64908)) ;
    dffr reg_ram_11__0 (.Q (ram_11__0), .QB (\$dummy [154]), .D (nx34630), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34631 (.Y (nx34630), .A0 (nx66026), .A1 (ram_11__0), .S0 (nx65182
             )) ;
    nand03 ix55058 (.Y (nx55057), .A0 (nx64870), .A1 (nx65368), .A2 (nx65140)) ;
    dffr reg_ram_10__0 (.Q (ram_10__0), .QB (\$dummy [155]), .D (nx34640), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34641 (.Y (nx34640), .A0 (nx66026), .A1 (ram_10__0), .S0 (nx65186
             )) ;
    nand03 ix55063 (.Y (nx55062), .A0 (nx64908), .A1 (nx65368), .A2 (nx65140)) ;
    aoi22 ix55066 (.Y (nx55065), .A0 (ram_12__0), .A1 (nx64946), .B0 (ram_13__0)
          , .B1 (nx64984)) ;
    dffr reg_ram_12__0 (.Q (ram_12__0), .QB (\$dummy [156]), .D (nx34620), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34621 (.Y (nx34620), .A0 (nx66026), .A1 (ram_12__0), .S0 (nx65190
             )) ;
    nand03 ix55070 (.Y (nx55069), .A0 (nx64946), .A1 (nx65368), .A2 (nx65140)) ;
    dffr reg_ram_13__0 (.Q (ram_13__0), .QB (\$dummy [157]), .D (nx34610), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34611 (.Y (nx34610), .A0 (nx66026), .A1 (ram_13__0), .S0 (nx65194
             )) ;
    nand03 ix55075 (.Y (nx55074), .A0 (nx64984), .A1 (nx65368), .A2 (nx65140)) ;
    aoi22 ix55078 (.Y (nx55077), .A0 (ram_15__0), .A1 (nx65022), .B0 (ram_14__0)
          , .B1 (nx65060)) ;
    dffr reg_ram_15__0 (.Q (ram_15__0), .QB (\$dummy [158]), .D (nx34590), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34591 (.Y (nx34590), .A0 (nx66026), .A1 (ram_15__0), .S0 (nx65198
             )) ;
    nand03 ix55082 (.Y (nx55081), .A0 (nx65022), .A1 (nx65370), .A2 (nx65142)) ;
    dffr reg_ram_14__0 (.Q (ram_14__0), .QB (\$dummy [159]), .D (nx34600), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34601 (.Y (nx34600), .A0 (nx66026), .A1 (ram_14__0), .S0 (nx65202
             )) ;
    nand03 ix55087 (.Y (nx55086), .A0 (nx65060), .A1 (nx65370), .A2 (nx65142)) ;
    oai21 ix55090 (.Y (nx55089), .A0 (nx1838), .A1 (nx1696), .B0 (nx65206)) ;
    nand04 ix1839 (.Y (nx1838), .A0 (nx55092), .A1 (nx55103), .A2 (nx55113), .A3 (
           nx55123)) ;
    aoi22 ix55093 (.Y (nx55092), .A0 (ram_96__0), .A1 (nx64490), .B0 (ram_97__0)
          , .B1 (nx64528)) ;
    dffr reg_ram_96__0 (.Q (ram_96__0), .QB (\$dummy [160]), .D (nx34580), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34581 (.Y (nx34580), .A0 (ram_96__0), .A1 (nx66026), .S0 (nx63784
             )) ;
    nand02 ix1555 (.Y (nx1554), .A0 (nx54554), .A1 (nx54282)) ;
    dffr reg_ram_97__0 (.Q (ram_97__0), .QB (\$dummy [161]), .D (nx34570), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34571 (.Y (nx34570), .A0 (ram_97__0), .A1 (nx66028), .S0 (nx63780
             )) ;
    aoi22 ix55104 (.Y (nx55103), .A0 (ram_99__0), .A1 (nx64566), .B0 (ram_98__0)
          , .B1 (nx64604)) ;
    dffr reg_ram_99__0 (.Q (ram_99__0), .QB (\$dummy [162]), .D (nx34550), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34551 (.Y (nx34550), .A0 (ram_99__0), .A1 (nx66028), .S0 (nx63772
             )) ;
    dffr reg_ram_98__0 (.Q (ram_98__0), .QB (\$dummy [163]), .D (nx34560), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34561 (.Y (nx34560), .A0 (ram_98__0), .A1 (nx66028), .S0 (nx63776
             )) ;
    aoi22 ix55114 (.Y (nx55113), .A0 (ram_100__0), .A1 (nx64642), .B0 (
          ram_101__0), .B1 (nx64680)) ;
    dffr reg_ram_100__0 (.Q (ram_100__0), .QB (\$dummy [164]), .D (nx34540), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34541 (.Y (nx34540), .A0 (ram_100__0), .A1 (nx66028), .S0 (
             nx63768)) ;
    dffr reg_ram_101__0 (.Q (ram_101__0), .QB (\$dummy [165]), .D (nx34530), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34531 (.Y (nx34530), .A0 (ram_101__0), .A1 (nx66028), .S0 (
             nx63764)) ;
    aoi22 ix55124 (.Y (nx55123), .A0 (ram_103__0), .A1 (nx64718), .B0 (
          ram_102__0), .B1 (nx64756)) ;
    dffr reg_ram_103__0 (.Q (ram_103__0), .QB (\$dummy [166]), .D (nx34510), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34511 (.Y (nx34510), .A0 (ram_103__0), .A1 (nx66028), .S0 (
             nx63756)) ;
    dffr reg_ram_102__0 (.Q (ram_102__0), .QB (\$dummy [167]), .D (nx34520), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34521 (.Y (nx34520), .A0 (ram_102__0), .A1 (nx66028), .S0 (
             nx63760)) ;
    nand04 ix1697 (.Y (nx1696), .A0 (nx55134), .A1 (nx55144), .A2 (nx55154), .A3 (
           nx55164)) ;
    aoi22 ix55135 (.Y (nx55134), .A0 (ram_104__0), .A1 (nx64794), .B0 (
          ram_105__0), .B1 (nx64832)) ;
    dffr reg_ram_104__0 (.Q (ram_104__0), .QB (\$dummy [168]), .D (nx34500), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34501 (.Y (nx34500), .A0 (ram_104__0), .A1 (nx66030), .S0 (
             nx63752)) ;
    dffr reg_ram_105__0 (.Q (ram_105__0), .QB (\$dummy [169]), .D (nx34490), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34491 (.Y (nx34490), .A0 (ram_105__0), .A1 (nx66030), .S0 (
             nx63748)) ;
    aoi22 ix55145 (.Y (nx55144), .A0 (ram_107__0), .A1 (nx64870), .B0 (
          ram_106__0), .B1 (nx64908)) ;
    dffr reg_ram_107__0 (.Q (ram_107__0), .QB (\$dummy [170]), .D (nx34470), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34471 (.Y (nx34470), .A0 (ram_107__0), .A1 (nx66030), .S0 (
             nx63740)) ;
    dffr reg_ram_106__0 (.Q (ram_106__0), .QB (\$dummy [171]), .D (nx34480), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34481 (.Y (nx34480), .A0 (ram_106__0), .A1 (nx66030), .S0 (
             nx63744)) ;
    aoi22 ix55155 (.Y (nx55154), .A0 (ram_108__0), .A1 (nx64946), .B0 (
          ram_109__0), .B1 (nx64984)) ;
    dffr reg_ram_108__0 (.Q (ram_108__0), .QB (\$dummy [172]), .D (nx34460), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34461 (.Y (nx34460), .A0 (ram_108__0), .A1 (nx66030), .S0 (
             nx63736)) ;
    dffr reg_ram_109__0 (.Q (ram_109__0), .QB (\$dummy [173]), .D (nx34450), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34451 (.Y (nx34450), .A0 (ram_109__0), .A1 (nx66030), .S0 (
             nx63732)) ;
    aoi22 ix55165 (.Y (nx55164), .A0 (ram_111__0), .A1 (nx65022), .B0 (
          ram_110__0), .B1 (nx65060)) ;
    dffr reg_ram_111__0 (.Q (ram_111__0), .QB (\$dummy [174]), .D (nx34430), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34431 (.Y (nx34430), .A0 (ram_111__0), .A1 (nx66030), .S0 (
             nx63724)) ;
    dffr reg_ram_110__0 (.Q (ram_110__0), .QB (\$dummy [175]), .D (nx34440), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34441 (.Y (nx34440), .A0 (ram_110__0), .A1 (nx66032), .S0 (
             nx63728)) ;
    oai21 ix55177 (.Y (nx55176), .A0 (nx1546), .A1 (nx1404), .B0 (nx65210)) ;
    nand04 ix1547 (.Y (nx1546), .A0 (nx55179), .A1 (nx55190), .A2 (nx55200), .A3 (
           nx55210)) ;
    aoi22 ix55180 (.Y (nx55179), .A0 (ram_112__0), .A1 (nx64490), .B0 (
          ram_113__0), .B1 (nx64528)) ;
    dffr reg_ram_112__0 (.Q (ram_112__0), .QB (\$dummy [176]), .D (nx34420), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34421 (.Y (nx34420), .A0 (ram_112__0), .A1 (nx66032), .S0 (
             nx63714)) ;
    nand03 ix1263 (.Y (nx1262), .A0 (nx54554), .A1 (address[4]), .A2 (nx65440)
           ) ;
    dffr reg_ram_113__0 (.Q (ram_113__0), .QB (\$dummy [177]), .D (nx34410), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34411 (.Y (nx34410), .A0 (ram_113__0), .A1 (nx66032), .S0 (
             nx63710)) ;
    aoi22 ix55191 (.Y (nx55190), .A0 (ram_115__0), .A1 (nx64566), .B0 (
          ram_114__0), .B1 (nx64604)) ;
    dffr reg_ram_115__0 (.Q (ram_115__0), .QB (\$dummy [178]), .D (nx34390), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34391 (.Y (nx34390), .A0 (ram_115__0), .A1 (nx66032), .S0 (
             nx63702)) ;
    dffr reg_ram_114__0 (.Q (ram_114__0), .QB (\$dummy [179]), .D (nx34400), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34401 (.Y (nx34400), .A0 (ram_114__0), .A1 (nx66032), .S0 (
             nx63706)) ;
    aoi22 ix55201 (.Y (nx55200), .A0 (ram_116__0), .A1 (nx64642), .B0 (
          ram_117__0), .B1 (nx64680)) ;
    dffr reg_ram_116__0 (.Q (ram_116__0), .QB (\$dummy [180]), .D (nx34380), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34381 (.Y (nx34380), .A0 (ram_116__0), .A1 (nx66032), .S0 (
             nx63698)) ;
    dffr reg_ram_117__0 (.Q (ram_117__0), .QB (\$dummy [181]), .D (nx34370), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34371 (.Y (nx34370), .A0 (ram_117__0), .A1 (nx66032), .S0 (
             nx63694)) ;
    aoi22 ix55211 (.Y (nx55210), .A0 (ram_119__0), .A1 (nx64718), .B0 (
          ram_118__0), .B1 (nx64756)) ;
    dffr reg_ram_119__0 (.Q (ram_119__0), .QB (\$dummy [182]), .D (nx34350), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34351 (.Y (nx34350), .A0 (ram_119__0), .A1 (nx66034), .S0 (
             nx63686)) ;
    dffr reg_ram_118__0 (.Q (ram_118__0), .QB (\$dummy [183]), .D (nx34360), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34361 (.Y (nx34360), .A0 (ram_118__0), .A1 (nx66034), .S0 (
             nx63690)) ;
    nand04 ix1405 (.Y (nx1404), .A0 (nx55221), .A1 (nx55231), .A2 (nx55241), .A3 (
           nx55251)) ;
    aoi22 ix55222 (.Y (nx55221), .A0 (ram_120__0), .A1 (nx64794), .B0 (
          ram_121__0), .B1 (nx64832)) ;
    dffr reg_ram_120__0 (.Q (ram_120__0), .QB (\$dummy [184]), .D (nx34340), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34341 (.Y (nx34340), .A0 (ram_120__0), .A1 (nx66034), .S0 (
             nx63682)) ;
    dffr reg_ram_121__0 (.Q (ram_121__0), .QB (\$dummy [185]), .D (nx34330), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34331 (.Y (nx34330), .A0 (ram_121__0), .A1 (nx66034), .S0 (
             nx63678)) ;
    aoi22 ix55232 (.Y (nx55231), .A0 (ram_123__0), .A1 (nx64870), .B0 (
          ram_122__0), .B1 (nx64908)) ;
    dffr reg_ram_123__0 (.Q (ram_123__0), .QB (\$dummy [186]), .D (nx34310), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34311 (.Y (nx34310), .A0 (ram_123__0), .A1 (nx66034), .S0 (
             nx63670)) ;
    dffr reg_ram_122__0 (.Q (ram_122__0), .QB (\$dummy [187]), .D (nx34320), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34321 (.Y (nx34320), .A0 (ram_122__0), .A1 (nx66034), .S0 (
             nx63674)) ;
    aoi22 ix55242 (.Y (nx55241), .A0 (ram_124__0), .A1 (nx64946), .B0 (
          ram_125__0), .B1 (nx64984)) ;
    dffr reg_ram_124__0 (.Q (ram_124__0), .QB (\$dummy [188]), .D (nx34300), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34301 (.Y (nx34300), .A0 (ram_124__0), .A1 (nx66034), .S0 (
             nx63666)) ;
    dffr reg_ram_125__0 (.Q (ram_125__0), .QB (\$dummy [189]), .D (nx34290), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34291 (.Y (nx34290), .A0 (ram_125__0), .A1 (nx66036), .S0 (
             nx63662)) ;
    aoi22 ix55252 (.Y (nx55251), .A0 (ram_127__0), .A1 (nx65022), .B0 (
          ram_126__0), .B1 (nx65060)) ;
    dffr reg_ram_127__0 (.Q (ram_127__0), .QB (\$dummy [190]), .D (nx34270), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34271 (.Y (nx34270), .A0 (ram_127__0), .A1 (nx66036), .S0 (
             nx63654)) ;
    dffr reg_ram_126__0 (.Q (ram_126__0), .QB (\$dummy [191]), .D (nx34280), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34281 (.Y (nx34280), .A0 (ram_126__0), .A1 (nx66036), .S0 (
             nx63658)) ;
    nand04 ix1257 (.Y (nx1256), .A0 (nx55264), .A1 (nx55355), .A2 (nx55442), .A3 (
           nx55529)) ;
    oai21 ix55265 (.Y (nx55264), .A0 (nx1246), .A1 (nx1104), .B0 (nx65214)) ;
    nand04 ix1247 (.Y (nx1246), .A0 (nx55267), .A1 (nx55282), .A2 (nx55292), .A3 (
           nx55302)) ;
    aoi22 ix55268 (.Y (nx55267), .A0 (ram_128__0), .A1 (nx64490), .B0 (
          ram_129__0), .B1 (nx64528)) ;
    dffr reg_ram_128__0 (.Q (ram_128__0), .QB (\$dummy [192]), .D (nx34260), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34261 (.Y (nx34260), .A0 (ram_128__0), .A1 (nx66036), .S0 (
             nx63644)) ;
    nand02 ix963 (.Y (nx962), .A0 (nx55273), .A1 (nx54464)) ;
    dffr reg_ram_129__0 (.Q (ram_129__0), .QB (\$dummy [193]), .D (nx34250), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34251 (.Y (nx34250), .A0 (ram_129__0), .A1 (nx66036), .S0 (
             nx63640)) ;
    aoi22 ix55283 (.Y (nx55282), .A0 (ram_131__0), .A1 (nx64566), .B0 (
          ram_130__0), .B1 (nx64604)) ;
    dffr reg_ram_131__0 (.Q (ram_131__0), .QB (\$dummy [194]), .D (nx34230), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34231 (.Y (nx34230), .A0 (ram_131__0), .A1 (nx66036), .S0 (
             nx63632)) ;
    dffr reg_ram_130__0 (.Q (ram_130__0), .QB (\$dummy [195]), .D (nx34240), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34241 (.Y (nx34240), .A0 (ram_130__0), .A1 (nx66036), .S0 (
             nx63636)) ;
    aoi22 ix55293 (.Y (nx55292), .A0 (ram_132__0), .A1 (nx64642), .B0 (
          ram_133__0), .B1 (nx64680)) ;
    dffr reg_ram_132__0 (.Q (ram_132__0), .QB (\$dummy [196]), .D (nx34220), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34221 (.Y (nx34220), .A0 (ram_132__0), .A1 (nx66038), .S0 (
             nx63628)) ;
    dffr reg_ram_133__0 (.Q (ram_133__0), .QB (\$dummy [197]), .D (nx34210), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34211 (.Y (nx34210), .A0 (ram_133__0), .A1 (nx66038), .S0 (
             nx63624)) ;
    aoi22 ix55303 (.Y (nx55302), .A0 (ram_135__0), .A1 (nx64718), .B0 (
          ram_134__0), .B1 (nx64756)) ;
    dffr reg_ram_135__0 (.Q (ram_135__0), .QB (\$dummy [198]), .D (nx34190), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34191 (.Y (nx34190), .A0 (ram_135__0), .A1 (nx66038), .S0 (
             nx63616)) ;
    dffr reg_ram_134__0 (.Q (ram_134__0), .QB (\$dummy [199]), .D (nx34200), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34201 (.Y (nx34200), .A0 (ram_134__0), .A1 (nx66038), .S0 (
             nx63620)) ;
    nand04 ix1105 (.Y (nx1104), .A0 (nx55313), .A1 (nx55323), .A2 (nx55333), .A3 (
           nx55343)) ;
    aoi22 ix55314 (.Y (nx55313), .A0 (ram_136__0), .A1 (nx64794), .B0 (
          ram_137__0), .B1 (nx64832)) ;
    dffr reg_ram_136__0 (.Q (ram_136__0), .QB (\$dummy [200]), .D (nx34180), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34181 (.Y (nx34180), .A0 (ram_136__0), .A1 (nx66038), .S0 (
             nx63612)) ;
    dffr reg_ram_137__0 (.Q (ram_137__0), .QB (\$dummy [201]), .D (nx34170), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34171 (.Y (nx34170), .A0 (ram_137__0), .A1 (nx66038), .S0 (
             nx63608)) ;
    aoi22 ix55324 (.Y (nx55323), .A0 (ram_139__0), .A1 (nx64870), .B0 (
          ram_138__0), .B1 (nx64908)) ;
    dffr reg_ram_139__0 (.Q (ram_139__0), .QB (\$dummy [202]), .D (nx34150), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34151 (.Y (nx34150), .A0 (ram_139__0), .A1 (nx66038), .S0 (
             nx63600)) ;
    dffr reg_ram_138__0 (.Q (ram_138__0), .QB (\$dummy [203]), .D (nx34160), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34161 (.Y (nx34160), .A0 (ram_138__0), .A1 (nx66040), .S0 (
             nx63604)) ;
    aoi22 ix55334 (.Y (nx55333), .A0 (ram_140__0), .A1 (nx64946), .B0 (
          ram_141__0), .B1 (nx64984)) ;
    dffr reg_ram_140__0 (.Q (ram_140__0), .QB (\$dummy [204]), .D (nx34140), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34141 (.Y (nx34140), .A0 (ram_140__0), .A1 (nx66040), .S0 (
             nx63596)) ;
    dffr reg_ram_141__0 (.Q (ram_141__0), .QB (\$dummy [205]), .D (nx34130), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34131 (.Y (nx34130), .A0 (ram_141__0), .A1 (nx66040), .S0 (
             nx63592)) ;
    aoi22 ix55344 (.Y (nx55343), .A0 (ram_143__0), .A1 (nx65022), .B0 (
          ram_142__0), .B1 (nx65060)) ;
    dffr reg_ram_143__0 (.Q (ram_143__0), .QB (\$dummy [206]), .D (nx34110), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34111 (.Y (nx34110), .A0 (ram_143__0), .A1 (nx66040), .S0 (
             nx63584)) ;
    dffr reg_ram_142__0 (.Q (ram_142__0), .QB (\$dummy [207]), .D (nx34120), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34121 (.Y (nx34120), .A0 (ram_142__0), .A1 (nx66040), .S0 (
             nx63588)) ;
    oai21 ix55356 (.Y (nx55355), .A0 (nx952), .A1 (nx810), .B0 (nx65218)) ;
    nand04 ix953 (.Y (nx952), .A0 (nx55358), .A1 (nx55369), .A2 (nx55379), .A3 (
           nx55389)) ;
    aoi22 ix55359 (.Y (nx55358), .A0 (ram_144__0), .A1 (nx64492), .B0 (
          ram_145__0), .B1 (nx64530)) ;
    dffr reg_ram_144__0 (.Q (ram_144__0), .QB (\$dummy [208]), .D (nx34100), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34101 (.Y (nx34100), .A0 (ram_144__0), .A1 (nx66040), .S0 (
             nx63574)) ;
    nand02 ix669 (.Y (nx668), .A0 (nx55273), .A1 (nx54373)) ;
    dffr reg_ram_145__0 (.Q (ram_145__0), .QB (\$dummy [209]), .D (nx34090), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34091 (.Y (nx34090), .A0 (ram_145__0), .A1 (nx66040), .S0 (
             nx63570)) ;
    aoi22 ix55370 (.Y (nx55369), .A0 (ram_147__0), .A1 (nx64568), .B0 (
          ram_146__0), .B1 (nx64606)) ;
    dffr reg_ram_147__0 (.Q (ram_147__0), .QB (\$dummy [210]), .D (nx34070), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34071 (.Y (nx34070), .A0 (ram_147__0), .A1 (nx66042), .S0 (
             nx63562)) ;
    dffr reg_ram_146__0 (.Q (ram_146__0), .QB (\$dummy [211]), .D (nx34080), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34081 (.Y (nx34080), .A0 (ram_146__0), .A1 (nx66042), .S0 (
             nx63566)) ;
    aoi22 ix55380 (.Y (nx55379), .A0 (ram_148__0), .A1 (nx64644), .B0 (
          ram_149__0), .B1 (nx64682)) ;
    dffr reg_ram_148__0 (.Q (ram_148__0), .QB (\$dummy [212]), .D (nx34060), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34061 (.Y (nx34060), .A0 (ram_148__0), .A1 (nx66042), .S0 (
             nx63558)) ;
    dffr reg_ram_149__0 (.Q (ram_149__0), .QB (\$dummy [213]), .D (nx34050), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34051 (.Y (nx34050), .A0 (ram_149__0), .A1 (nx66042), .S0 (
             nx63554)) ;
    aoi22 ix55390 (.Y (nx55389), .A0 (ram_151__0), .A1 (nx64720), .B0 (
          ram_150__0), .B1 (nx64758)) ;
    dffr reg_ram_151__0 (.Q (ram_151__0), .QB (\$dummy [214]), .D (nx34030), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34031 (.Y (nx34030), .A0 (ram_151__0), .A1 (nx66042), .S0 (
             nx63546)) ;
    dffr reg_ram_150__0 (.Q (ram_150__0), .QB (\$dummy [215]), .D (nx34040), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34041 (.Y (nx34040), .A0 (ram_150__0), .A1 (nx66042), .S0 (
             nx63550)) ;
    nand04 ix811 (.Y (nx810), .A0 (nx55400), .A1 (nx55410), .A2 (nx55420), .A3 (
           nx55430)) ;
    aoi22 ix55401 (.Y (nx55400), .A0 (ram_152__0), .A1 (nx64796), .B0 (
          ram_153__0), .B1 (nx64834)) ;
    dffr reg_ram_152__0 (.Q (ram_152__0), .QB (\$dummy [216]), .D (nx34020), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34021 (.Y (nx34020), .A0 (ram_152__0), .A1 (nx66042), .S0 (
             nx63542)) ;
    dffr reg_ram_153__0 (.Q (ram_153__0), .QB (\$dummy [217]), .D (nx34010), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34011 (.Y (nx34010), .A0 (ram_153__0), .A1 (nx66044), .S0 (
             nx63538)) ;
    aoi22 ix55411 (.Y (nx55410), .A0 (ram_155__0), .A1 (nx64872), .B0 (
          ram_154__0), .B1 (nx64910)) ;
    dffr reg_ram_155__0 (.Q (ram_155__0), .QB (\$dummy [218]), .D (nx33990), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33991 (.Y (nx33990), .A0 (ram_155__0), .A1 (nx66044), .S0 (
             nx63530)) ;
    dffr reg_ram_154__0 (.Q (ram_154__0), .QB (\$dummy [219]), .D (nx34000), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix34001 (.Y (nx34000), .A0 (ram_154__0), .A1 (nx66044), .S0 (
             nx63534)) ;
    aoi22 ix55421 (.Y (nx55420), .A0 (ram_156__0), .A1 (nx64948), .B0 (
          ram_157__0), .B1 (nx64986)) ;
    dffr reg_ram_156__0 (.Q (ram_156__0), .QB (\$dummy [220]), .D (nx33980), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33981 (.Y (nx33980), .A0 (ram_156__0), .A1 (nx66044), .S0 (
             nx63526)) ;
    dffr reg_ram_157__0 (.Q (ram_157__0), .QB (\$dummy [221]), .D (nx33970), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33971 (.Y (nx33970), .A0 (ram_157__0), .A1 (nx66044), .S0 (
             nx63522)) ;
    aoi22 ix55431 (.Y (nx55430), .A0 (ram_159__0), .A1 (nx65024), .B0 (
          ram_158__0), .B1 (nx65062)) ;
    dffr reg_ram_159__0 (.Q (ram_159__0), .QB (\$dummy [222]), .D (nx33950), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33951 (.Y (nx33950), .A0 (ram_159__0), .A1 (nx66044), .S0 (
             nx63514)) ;
    dffr reg_ram_158__0 (.Q (ram_158__0), .QB (\$dummy [223]), .D (nx33960), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33961 (.Y (nx33960), .A0 (ram_158__0), .A1 (nx66044), .S0 (
             nx63518)) ;
    oai21 ix55443 (.Y (nx55442), .A0 (nx654), .A1 (nx512), .B0 (nx65222)) ;
    nand04 ix655 (.Y (nx654), .A0 (nx55445), .A1 (nx55456), .A2 (nx55466), .A3 (
           nx55476)) ;
    aoi22 ix55446 (.Y (nx55445), .A0 (ram_160__0), .A1 (nx64492), .B0 (
          ram_161__0), .B1 (nx64530)) ;
    dffr reg_ram_160__0 (.Q (ram_160__0), .QB (\$dummy [224]), .D (nx33940), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33941 (.Y (nx33940), .A0 (ram_160__0), .A1 (nx66046), .S0 (
             nx63504)) ;
    nand02 ix371 (.Y (nx370), .A0 (nx55273), .A1 (nx54282)) ;
    dffr reg_ram_161__0 (.Q (ram_161__0), .QB (\$dummy [225]), .D (nx33930), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33931 (.Y (nx33930), .A0 (ram_161__0), .A1 (nx66046), .S0 (
             nx63500)) ;
    aoi22 ix55457 (.Y (nx55456), .A0 (ram_163__0), .A1 (nx64568), .B0 (
          ram_162__0), .B1 (nx64606)) ;
    dffr reg_ram_163__0 (.Q (ram_163__0), .QB (\$dummy [226]), .D (nx33910), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33911 (.Y (nx33910), .A0 (ram_163__0), .A1 (nx66046), .S0 (
             nx63492)) ;
    dffr reg_ram_162__0 (.Q (ram_162__0), .QB (\$dummy [227]), .D (nx33920), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33921 (.Y (nx33920), .A0 (ram_162__0), .A1 (nx66046), .S0 (
             nx63496)) ;
    aoi22 ix55467 (.Y (nx55466), .A0 (ram_164__0), .A1 (nx64644), .B0 (
          ram_165__0), .B1 (nx64682)) ;
    dffr reg_ram_164__0 (.Q (ram_164__0), .QB (\$dummy [228]), .D (nx33900), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33901 (.Y (nx33900), .A0 (ram_164__0), .A1 (nx66046), .S0 (
             nx63488)) ;
    dffr reg_ram_165__0 (.Q (ram_165__0), .QB (\$dummy [229]), .D (nx33890), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33891 (.Y (nx33890), .A0 (ram_165__0), .A1 (nx66046), .S0 (
             nx63484)) ;
    aoi22 ix55477 (.Y (nx55476), .A0 (ram_167__0), .A1 (nx64720), .B0 (
          ram_166__0), .B1 (nx64758)) ;
    dffr reg_ram_167__0 (.Q (ram_167__0), .QB (\$dummy [230]), .D (nx33870), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33871 (.Y (nx33870), .A0 (ram_167__0), .A1 (nx66046), .S0 (
             nx63476)) ;
    dffr reg_ram_166__0 (.Q (ram_166__0), .QB (\$dummy [231]), .D (nx33880), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33881 (.Y (nx33880), .A0 (ram_166__0), .A1 (nx66048), .S0 (
             nx63480)) ;
    nand04 ix513 (.Y (nx512), .A0 (nx55487), .A1 (nx55497), .A2 (nx55507), .A3 (
           nx55517)) ;
    aoi22 ix55488 (.Y (nx55487), .A0 (ram_168__0), .A1 (nx64796), .B0 (
          ram_169__0), .B1 (nx64834)) ;
    dffr reg_ram_168__0 (.Q (ram_168__0), .QB (\$dummy [232]), .D (nx33860), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33861 (.Y (nx33860), .A0 (ram_168__0), .A1 (nx66048), .S0 (
             nx63472)) ;
    dffr reg_ram_169__0 (.Q (ram_169__0), .QB (\$dummy [233]), .D (nx33850), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33851 (.Y (nx33850), .A0 (ram_169__0), .A1 (nx66048), .S0 (
             nx63468)) ;
    aoi22 ix55498 (.Y (nx55497), .A0 (ram_171__0), .A1 (nx64872), .B0 (
          ram_170__0), .B1 (nx64910)) ;
    dffr reg_ram_171__0 (.Q (ram_171__0), .QB (\$dummy [234]), .D (nx33830), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33831 (.Y (nx33830), .A0 (ram_171__0), .A1 (nx66048), .S0 (
             nx63460)) ;
    dffr reg_ram_170__0 (.Q (ram_170__0), .QB (\$dummy [235]), .D (nx33840), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33841 (.Y (nx33840), .A0 (ram_170__0), .A1 (nx66048), .S0 (
             nx63464)) ;
    aoi22 ix55508 (.Y (nx55507), .A0 (ram_172__0), .A1 (nx64948), .B0 (
          ram_173__0), .B1 (nx64986)) ;
    dffr reg_ram_172__0 (.Q (ram_172__0), .QB (\$dummy [236]), .D (nx33820), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33821 (.Y (nx33820), .A0 (ram_172__0), .A1 (nx66048), .S0 (
             nx63456)) ;
    dffr reg_ram_173__0 (.Q (ram_173__0), .QB (\$dummy [237]), .D (nx33810), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33811 (.Y (nx33810), .A0 (ram_173__0), .A1 (nx66048), .S0 (
             nx63452)) ;
    aoi22 ix55518 (.Y (nx55517), .A0 (ram_175__0), .A1 (nx65024), .B0 (
          ram_174__0), .B1 (nx65062)) ;
    dffr reg_ram_175__0 (.Q (ram_175__0), .QB (\$dummy [238]), .D (nx33790), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33791 (.Y (nx33790), .A0 (ram_175__0), .A1 (nx66050), .S0 (
             nx63444)) ;
    dffr reg_ram_174__0 (.Q (ram_174__0), .QB (\$dummy [239]), .D (nx33800), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33801 (.Y (nx33800), .A0 (ram_174__0), .A1 (nx66050), .S0 (
             nx63448)) ;
    oai21 ix55530 (.Y (nx55529), .A0 (nx358), .A1 (nx194), .B0 (nx65226)) ;
    nand04 ix359 (.Y (nx358), .A0 (nx55532), .A1 (nx55543), .A2 (nx55553), .A3 (
           nx55563)) ;
    aoi22 ix55533 (.Y (nx55532), .A0 (ram_176__0), .A1 (nx64492), .B0 (
          ram_177__0), .B1 (nx64530)) ;
    dffr reg_ram_176__0 (.Q (ram_176__0), .QB (\$dummy [240]), .D (nx33780), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33781 (.Y (nx33780), .A0 (ram_176__0), .A1 (nx66050), .S0 (
             nx63434)) ;
    nand03 ix11 (.Y (nx10), .A0 (nx55273), .A1 (address[4]), .A2 (nx65440)) ;
    dffr reg_ram_177__0 (.Q (ram_177__0), .QB (\$dummy [241]), .D (nx33770), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33771 (.Y (nx33770), .A0 (ram_177__0), .A1 (nx66050), .S0 (
             nx63424)) ;
    aoi22 ix55544 (.Y (nx55543), .A0 (ram_179__0), .A1 (nx64568), .B0 (
          ram_178__0), .B1 (nx64606)) ;
    dffr reg_ram_179__0 (.Q (ram_179__0), .QB (\$dummy [242]), .D (nx33750), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33751 (.Y (nx33750), .A0 (ram_179__0), .A1 (nx66050), .S0 (
             nx63404)) ;
    dffr reg_ram_178__0 (.Q (ram_178__0), .QB (\$dummy [243]), .D (nx33760), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33761 (.Y (nx33760), .A0 (ram_178__0), .A1 (nx66050), .S0 (
             nx63414)) ;
    aoi22 ix55554 (.Y (nx55553), .A0 (ram_180__0), .A1 (nx64644), .B0 (
          ram_181__0), .B1 (nx64682)) ;
    dffr reg_ram_180__0 (.Q (ram_180__0), .QB (\$dummy [244]), .D (nx33740), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33741 (.Y (nx33740), .A0 (ram_180__0), .A1 (nx66050), .S0 (
             nx63394)) ;
    dffr reg_ram_181__0 (.Q (ram_181__0), .QB (\$dummy [245]), .D (nx33730), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33731 (.Y (nx33730), .A0 (ram_181__0), .A1 (nx66052), .S0 (
             nx63384)) ;
    aoi22 ix55564 (.Y (nx55563), .A0 (ram_183__0), .A1 (nx64720), .B0 (
          ram_182__0), .B1 (nx64758)) ;
    dffr reg_ram_183__0 (.Q (ram_183__0), .QB (\$dummy [246]), .D (nx33710), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33711 (.Y (nx33710), .A0 (ram_183__0), .A1 (nx66052), .S0 (
             nx63364)) ;
    dffr reg_ram_182__0 (.Q (ram_182__0), .QB (\$dummy [247]), .D (nx33720), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33721 (.Y (nx33720), .A0 (ram_182__0), .A1 (nx66052), .S0 (
             nx63374)) ;
    nand04 ix195 (.Y (nx194), .A0 (nx55574), .A1 (nx55584), .A2 (nx55594), .A3 (
           nx55604)) ;
    aoi22 ix55575 (.Y (nx55574), .A0 (ram_184__0), .A1 (nx64796), .B0 (
          ram_185__0), .B1 (nx64834)) ;
    dffr reg_ram_184__0 (.Q (ram_184__0), .QB (\$dummy [248]), .D (nx33700), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33701 (.Y (nx33700), .A0 (ram_184__0), .A1 (nx66052), .S0 (
             nx63354)) ;
    dffr reg_ram_185__0 (.Q (ram_185__0), .QB (\$dummy [249]), .D (nx33690), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33691 (.Y (nx33690), .A0 (ram_185__0), .A1 (nx66052), .S0 (
             nx63344)) ;
    aoi22 ix55585 (.Y (nx55584), .A0 (ram_187__0), .A1 (nx64872), .B0 (
          ram_186__0), .B1 (nx64910)) ;
    dffr reg_ram_187__0 (.Q (ram_187__0), .QB (\$dummy [250]), .D (nx33670), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33671 (.Y (nx33670), .A0 (ram_187__0), .A1 (nx66052), .S0 (
             nx63324)) ;
    dffr reg_ram_186__0 (.Q (ram_186__0), .QB (\$dummy [251]), .D (nx33680), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33681 (.Y (nx33680), .A0 (ram_186__0), .A1 (nx66052), .S0 (
             nx63334)) ;
    aoi22 ix55595 (.Y (nx55594), .A0 (ram_188__0), .A1 (nx64948), .B0 (
          ram_189__0), .B1 (nx64986)) ;
    dffr reg_ram_188__0 (.Q (ram_188__0), .QB (\$dummy [252]), .D (nx33660), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33661 (.Y (nx33660), .A0 (ram_188__0), .A1 (nx66054), .S0 (
             nx63314)) ;
    dffr reg_ram_189__0 (.Q (ram_189__0), .QB (\$dummy [253]), .D (nx33650), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33651 (.Y (nx33650), .A0 (ram_189__0), .A1 (nx66054), .S0 (
             nx63304)) ;
    aoi22 ix55605 (.Y (nx55604), .A0 (ram_191__0), .A1 (nx65024), .B0 (
          ram_190__0), .B1 (nx65062)) ;
    dffr reg_ram_191__0 (.Q (ram_191__0), .QB (\$dummy [254]), .D (nx33630), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33631 (.Y (nx33630), .A0 (ram_191__0), .A1 (nx66054), .S0 (
             nx63284)) ;
    dffr reg_ram_190__0 (.Q (ram_190__0), .QB (\$dummy [255]), .D (nx33640), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix33641 (.Y (nx33640), .A0 (ram_190__0), .A1 (nx66054), .S0 (
             nx63294)) ;
    or04 ix7419 (.Y (dataout[1]), .A0 (nx7414), .A1 (nx6760), .A2 (nx6104), .A3 (
         nx5450)) ;
    nand04 ix7415 (.Y (nx7414), .A0 (nx55618), .A1 (nx55686), .A2 (nx55754), .A3 (
           nx55822)) ;
    oai21 ix55619 (.Y (nx55618), .A0 (nx7404), .A1 (nx7326), .B0 (nx65096)) ;
    nand04 ix7405 (.Y (nx7404), .A0 (nx55621), .A1 (nx55629), .A2 (nx55637), .A3 (
           nx55645)) ;
    aoi22 ix55622 (.Y (nx55621), .A0 (ram_240__1), .A1 (nx64492), .B0 (
          ram_241__1), .B1 (nx64530)) ;
    dffr reg_ram_240__1 (.Q (ram_240__1), .QB (\$dummy [256]), .D (nx38740), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38741 (.Y (nx38740), .A0 (ram_240__1), .A1 (nx65906), .S0 (
             nx64414)) ;
    dffr reg_ram_241__1 (.Q (ram_241__1), .QB (\$dummy [257]), .D (nx38730), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38731 (.Y (nx38730), .A0 (ram_241__1), .A1 (nx65906), .S0 (
             nx64410)) ;
    aoi22 ix55630 (.Y (nx55629), .A0 (ram_243__1), .A1 (nx64568), .B0 (
          ram_242__1), .B1 (nx64606)) ;
    dffr reg_ram_243__1 (.Q (ram_243__1), .QB (\$dummy [258]), .D (nx38710), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38711 (.Y (nx38710), .A0 (ram_243__1), .A1 (nx65906), .S0 (
             nx64402)) ;
    dffr reg_ram_242__1 (.Q (ram_242__1), .QB (\$dummy [259]), .D (nx38720), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38721 (.Y (nx38720), .A0 (ram_242__1), .A1 (nx65906), .S0 (
             nx64406)) ;
    aoi22 ix55638 (.Y (nx55637), .A0 (ram_244__1), .A1 (nx64644), .B0 (
          ram_245__1), .B1 (nx64682)) ;
    dffr reg_ram_244__1 (.Q (ram_244__1), .QB (\$dummy [260]), .D (nx38700), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38701 (.Y (nx38700), .A0 (ram_244__1), .A1 (nx65906), .S0 (
             nx64398)) ;
    dffr reg_ram_245__1 (.Q (ram_245__1), .QB (\$dummy [261]), .D (nx38690), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38691 (.Y (nx38690), .A0 (ram_245__1), .A1 (nx65906), .S0 (
             nx64394)) ;
    aoi22 ix55646 (.Y (nx55645), .A0 (ram_247__1), .A1 (nx64720), .B0 (
          ram_246__1), .B1 (nx64758)) ;
    dffr reg_ram_247__1 (.Q (ram_247__1), .QB (\$dummy [262]), .D (nx38670), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38671 (.Y (nx38670), .A0 (ram_247__1), .A1 (nx65906), .S0 (
             nx64386)) ;
    dffr reg_ram_246__1 (.Q (ram_246__1), .QB (\$dummy [263]), .D (nx38680), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38681 (.Y (nx38680), .A0 (ram_246__1), .A1 (nx65908), .S0 (
             nx64390)) ;
    nand04 ix7327 (.Y (nx7326), .A0 (nx55654), .A1 (nx55662), .A2 (nx55670), .A3 (
           nx55678)) ;
    aoi22 ix55655 (.Y (nx55654), .A0 (ram_248__1), .A1 (nx64796), .B0 (
          ram_249__1), .B1 (nx64834)) ;
    dffr reg_ram_248__1 (.Q (ram_248__1), .QB (\$dummy [264]), .D (nx38660), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38661 (.Y (nx38660), .A0 (ram_248__1), .A1 (nx65908), .S0 (
             nx64382)) ;
    dffr reg_ram_249__1 (.Q (ram_249__1), .QB (\$dummy [265]), .D (nx38650), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38651 (.Y (nx38650), .A0 (ram_249__1), .A1 (nx65908), .S0 (
             nx64378)) ;
    aoi22 ix55663 (.Y (nx55662), .A0 (ram_251__1), .A1 (nx64872), .B0 (
          ram_250__1), .B1 (nx64910)) ;
    dffr reg_ram_251__1 (.Q (ram_251__1), .QB (\$dummy [266]), .D (nx38630), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38631 (.Y (nx38630), .A0 (ram_251__1), .A1 (nx65908), .S0 (
             nx64370)) ;
    dffr reg_ram_250__1 (.Q (ram_250__1), .QB (\$dummy [267]), .D (nx38640), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38641 (.Y (nx38640), .A0 (ram_250__1), .A1 (nx65908), .S0 (
             nx64374)) ;
    aoi22 ix55671 (.Y (nx55670), .A0 (ram_252__1), .A1 (nx64948), .B0 (
          ram_253__1), .B1 (nx64986)) ;
    dffr reg_ram_252__1 (.Q (ram_252__1), .QB (\$dummy [268]), .D (nx38620), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38621 (.Y (nx38620), .A0 (ram_252__1), .A1 (nx65908), .S0 (
             nx64366)) ;
    dffr reg_ram_253__1 (.Q (ram_253__1), .QB (\$dummy [269]), .D (nx38610), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38611 (.Y (nx38610), .A0 (ram_253__1), .A1 (nx65908), .S0 (
             nx64362)) ;
    aoi22 ix55679 (.Y (nx55678), .A0 (ram_255__1), .A1 (nx65024), .B0 (
          ram_254__1), .B1 (nx65062)) ;
    dffr reg_ram_255__1 (.Q (ram_255__1), .QB (\$dummy [270]), .D (nx38590), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38591 (.Y (nx38590), .A0 (ram_255__1), .A1 (nx65910), .S0 (
             nx64354)) ;
    dffr reg_ram_254__1 (.Q (ram_254__1), .QB (\$dummy [271]), .D (nx38600), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38601 (.Y (nx38600), .A0 (ram_254__1), .A1 (nx65910), .S0 (
             nx64358)) ;
    oai21 ix55687 (.Y (nx55686), .A0 (nx7242), .A1 (nx7164), .B0 (nx65100)) ;
    nand04 ix7243 (.Y (nx7242), .A0 (nx55689), .A1 (nx55697), .A2 (nx55705), .A3 (
           nx55713)) ;
    aoi22 ix55690 (.Y (nx55689), .A0 (ram_224__1), .A1 (nx64492), .B0 (
          ram_225__1), .B1 (nx64530)) ;
    dffr reg_ram_224__1 (.Q (ram_224__1), .QB (\$dummy [272]), .D (nx38580), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38581 (.Y (nx38580), .A0 (ram_224__1), .A1 (nx65910), .S0 (
             nx64344)) ;
    dffr reg_ram_225__1 (.Q (ram_225__1), .QB (\$dummy [273]), .D (nx38570), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38571 (.Y (nx38570), .A0 (ram_225__1), .A1 (nx65910), .S0 (
             nx64340)) ;
    aoi22 ix55698 (.Y (nx55697), .A0 (ram_227__1), .A1 (nx64568), .B0 (
          ram_226__1), .B1 (nx64606)) ;
    dffr reg_ram_227__1 (.Q (ram_227__1), .QB (\$dummy [274]), .D (nx38550), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38551 (.Y (nx38550), .A0 (ram_227__1), .A1 (nx65910), .S0 (
             nx64332)) ;
    dffr reg_ram_226__1 (.Q (ram_226__1), .QB (\$dummy [275]), .D (nx38560), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38561 (.Y (nx38560), .A0 (ram_226__1), .A1 (nx65910), .S0 (
             nx64336)) ;
    aoi22 ix55706 (.Y (nx55705), .A0 (ram_228__1), .A1 (nx64644), .B0 (
          ram_229__1), .B1 (nx64682)) ;
    dffr reg_ram_228__1 (.Q (ram_228__1), .QB (\$dummy [276]), .D (nx38540), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38541 (.Y (nx38540), .A0 (ram_228__1), .A1 (nx65910), .S0 (
             nx64328)) ;
    dffr reg_ram_229__1 (.Q (ram_229__1), .QB (\$dummy [277]), .D (nx38530), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38531 (.Y (nx38530), .A0 (ram_229__1), .A1 (nx65912), .S0 (
             nx64324)) ;
    aoi22 ix55714 (.Y (nx55713), .A0 (ram_231__1), .A1 (nx64720), .B0 (
          ram_230__1), .B1 (nx64758)) ;
    dffr reg_ram_231__1 (.Q (ram_231__1), .QB (\$dummy [278]), .D (nx38510), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38511 (.Y (nx38510), .A0 (ram_231__1), .A1 (nx65912), .S0 (
             nx64316)) ;
    dffr reg_ram_230__1 (.Q (ram_230__1), .QB (\$dummy [279]), .D (nx38520), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38521 (.Y (nx38520), .A0 (ram_230__1), .A1 (nx65912), .S0 (
             nx64320)) ;
    nand04 ix7165 (.Y (nx7164), .A0 (nx55722), .A1 (nx55730), .A2 (nx55738), .A3 (
           nx55746)) ;
    aoi22 ix55723 (.Y (nx55722), .A0 (ram_232__1), .A1 (nx64796), .B0 (
          ram_233__1), .B1 (nx64834)) ;
    dffr reg_ram_232__1 (.Q (ram_232__1), .QB (\$dummy [280]), .D (nx38500), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38501 (.Y (nx38500), .A0 (ram_232__1), .A1 (nx65912), .S0 (
             nx64312)) ;
    dffr reg_ram_233__1 (.Q (ram_233__1), .QB (\$dummy [281]), .D (nx38490), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38491 (.Y (nx38490), .A0 (ram_233__1), .A1 (nx65912), .S0 (
             nx64308)) ;
    aoi22 ix55731 (.Y (nx55730), .A0 (ram_235__1), .A1 (nx64872), .B0 (
          ram_234__1), .B1 (nx64910)) ;
    dffr reg_ram_235__1 (.Q (ram_235__1), .QB (\$dummy [282]), .D (nx38470), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38471 (.Y (nx38470), .A0 (ram_235__1), .A1 (nx65912), .S0 (
             nx64300)) ;
    dffr reg_ram_234__1 (.Q (ram_234__1), .QB (\$dummy [283]), .D (nx38480), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38481 (.Y (nx38480), .A0 (ram_234__1), .A1 (nx65912), .S0 (
             nx64304)) ;
    aoi22 ix55739 (.Y (nx55738), .A0 (ram_236__1), .A1 (nx64948), .B0 (
          ram_237__1), .B1 (nx64986)) ;
    dffr reg_ram_236__1 (.Q (ram_236__1), .QB (\$dummy [284]), .D (nx38460), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38461 (.Y (nx38460), .A0 (ram_236__1), .A1 (nx65914), .S0 (
             nx64296)) ;
    dffr reg_ram_237__1 (.Q (ram_237__1), .QB (\$dummy [285]), .D (nx38450), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38451 (.Y (nx38450), .A0 (ram_237__1), .A1 (nx65914), .S0 (
             nx64292)) ;
    aoi22 ix55747 (.Y (nx55746), .A0 (ram_239__1), .A1 (nx65024), .B0 (
          ram_238__1), .B1 (nx65062)) ;
    dffr reg_ram_239__1 (.Q (ram_239__1), .QB (\$dummy [286]), .D (nx38430), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38431 (.Y (nx38430), .A0 (ram_239__1), .A1 (nx65914), .S0 (
             nx64284)) ;
    dffr reg_ram_238__1 (.Q (ram_238__1), .QB (\$dummy [287]), .D (nx38440), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38441 (.Y (nx38440), .A0 (ram_238__1), .A1 (nx65914), .S0 (
             nx64288)) ;
    oai21 ix55755 (.Y (nx55754), .A0 (nx7078), .A1 (nx7000), .B0 (nx65104)) ;
    nand04 ix7079 (.Y (nx7078), .A0 (nx55757), .A1 (nx55765), .A2 (nx55773), .A3 (
           nx55781)) ;
    aoi22 ix55758 (.Y (nx55757), .A0 (ram_208__1), .A1 (nx64492), .B0 (
          ram_209__1), .B1 (nx64530)) ;
    dffr reg_ram_208__1 (.Q (ram_208__1), .QB (\$dummy [288]), .D (nx38420), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38421 (.Y (nx38420), .A0 (ram_208__1), .A1 (nx65914), .S0 (
             nx64274)) ;
    dffr reg_ram_209__1 (.Q (ram_209__1), .QB (\$dummy [289]), .D (nx38410), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38411 (.Y (nx38410), .A0 (ram_209__1), .A1 (nx65914), .S0 (
             nx64270)) ;
    aoi22 ix55766 (.Y (nx55765), .A0 (ram_211__1), .A1 (nx64568), .B0 (
          ram_210__1), .B1 (nx64606)) ;
    dffr reg_ram_211__1 (.Q (ram_211__1), .QB (\$dummy [290]), .D (nx38390), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38391 (.Y (nx38390), .A0 (ram_211__1), .A1 (nx65914), .S0 (
             nx64262)) ;
    dffr reg_ram_210__1 (.Q (ram_210__1), .QB (\$dummy [291]), .D (nx38400), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38401 (.Y (nx38400), .A0 (ram_210__1), .A1 (nx65916), .S0 (
             nx64266)) ;
    aoi22 ix55774 (.Y (nx55773), .A0 (ram_212__1), .A1 (nx64644), .B0 (
          ram_213__1), .B1 (nx64682)) ;
    dffr reg_ram_212__1 (.Q (ram_212__1), .QB (\$dummy [292]), .D (nx38380), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38381 (.Y (nx38380), .A0 (ram_212__1), .A1 (nx65916), .S0 (
             nx64258)) ;
    dffr reg_ram_213__1 (.Q (ram_213__1), .QB (\$dummy [293]), .D (nx38370), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38371 (.Y (nx38370), .A0 (ram_213__1), .A1 (nx65916), .S0 (
             nx64254)) ;
    aoi22 ix55782 (.Y (nx55781), .A0 (ram_215__1), .A1 (nx64720), .B0 (
          ram_214__1), .B1 (nx64758)) ;
    dffr reg_ram_215__1 (.Q (ram_215__1), .QB (\$dummy [294]), .D (nx38350), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38351 (.Y (nx38350), .A0 (ram_215__1), .A1 (nx65916), .S0 (
             nx64246)) ;
    dffr reg_ram_214__1 (.Q (ram_214__1), .QB (\$dummy [295]), .D (nx38360), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38361 (.Y (nx38360), .A0 (ram_214__1), .A1 (nx65916), .S0 (
             nx64250)) ;
    nand04 ix7001 (.Y (nx7000), .A0 (nx55790), .A1 (nx55798), .A2 (nx55806), .A3 (
           nx55814)) ;
    aoi22 ix55791 (.Y (nx55790), .A0 (ram_216__1), .A1 (nx64796), .B0 (
          ram_217__1), .B1 (nx64834)) ;
    dffr reg_ram_216__1 (.Q (ram_216__1), .QB (\$dummy [296]), .D (nx38340), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38341 (.Y (nx38340), .A0 (ram_216__1), .A1 (nx65916), .S0 (
             nx64242)) ;
    dffr reg_ram_217__1 (.Q (ram_217__1), .QB (\$dummy [297]), .D (nx38330), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38331 (.Y (nx38330), .A0 (ram_217__1), .A1 (nx65916), .S0 (
             nx64238)) ;
    aoi22 ix55799 (.Y (nx55798), .A0 (ram_219__1), .A1 (nx64872), .B0 (
          ram_218__1), .B1 (nx64910)) ;
    dffr reg_ram_219__1 (.Q (ram_219__1), .QB (\$dummy [298]), .D (nx38310), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38311 (.Y (nx38310), .A0 (ram_219__1), .A1 (nx65918), .S0 (
             nx64230)) ;
    dffr reg_ram_218__1 (.Q (ram_218__1), .QB (\$dummy [299]), .D (nx38320), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38321 (.Y (nx38320), .A0 (ram_218__1), .A1 (nx65918), .S0 (
             nx64234)) ;
    aoi22 ix55807 (.Y (nx55806), .A0 (ram_220__1), .A1 (nx64948), .B0 (
          ram_221__1), .B1 (nx64986)) ;
    dffr reg_ram_220__1 (.Q (ram_220__1), .QB (\$dummy [300]), .D (nx38300), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38301 (.Y (nx38300), .A0 (ram_220__1), .A1 (nx65918), .S0 (
             nx64226)) ;
    dffr reg_ram_221__1 (.Q (ram_221__1), .QB (\$dummy [301]), .D (nx38290), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38291 (.Y (nx38290), .A0 (ram_221__1), .A1 (nx65918), .S0 (
             nx64222)) ;
    aoi22 ix55815 (.Y (nx55814), .A0 (ram_223__1), .A1 (nx65024), .B0 (
          ram_222__1), .B1 (nx65062)) ;
    dffr reg_ram_223__1 (.Q (ram_223__1), .QB (\$dummy [302]), .D (nx38270), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38271 (.Y (nx38270), .A0 (ram_223__1), .A1 (nx65918), .S0 (
             nx64214)) ;
    dffr reg_ram_222__1 (.Q (ram_222__1), .QB (\$dummy [303]), .D (nx38280), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38281 (.Y (nx38280), .A0 (ram_222__1), .A1 (nx65918), .S0 (
             nx64218)) ;
    oai21 ix55823 (.Y (nx55822), .A0 (nx6916), .A1 (nx6838), .B0 (nx65108)) ;
    nand04 ix6917 (.Y (nx6916), .A0 (nx55825), .A1 (nx55833), .A2 (nx55841), .A3 (
           nx55849)) ;
    aoi22 ix55826 (.Y (nx55825), .A0 (ram_192__1), .A1 (nx64492), .B0 (
          ram_193__1), .B1 (nx64530)) ;
    dffr reg_ram_192__1 (.Q (ram_192__1), .QB (\$dummy [304]), .D (nx38260), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38261 (.Y (nx38260), .A0 (ram_192__1), .A1 (nx65918), .S0 (
             nx64204)) ;
    dffr reg_ram_193__1 (.Q (ram_193__1), .QB (\$dummy [305]), .D (nx38250), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38251 (.Y (nx38250), .A0 (ram_193__1), .A1 (nx65920), .S0 (
             nx64200)) ;
    aoi22 ix55834 (.Y (nx55833), .A0 (ram_195__1), .A1 (nx64568), .B0 (
          ram_194__1), .B1 (nx64606)) ;
    dffr reg_ram_195__1 (.Q (ram_195__1), .QB (\$dummy [306]), .D (nx38230), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38231 (.Y (nx38230), .A0 (ram_195__1), .A1 (nx65920), .S0 (
             nx64192)) ;
    dffr reg_ram_194__1 (.Q (ram_194__1), .QB (\$dummy [307]), .D (nx38240), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38241 (.Y (nx38240), .A0 (ram_194__1), .A1 (nx65920), .S0 (
             nx64196)) ;
    aoi22 ix55842 (.Y (nx55841), .A0 (ram_196__1), .A1 (nx64644), .B0 (
          ram_197__1), .B1 (nx64682)) ;
    dffr reg_ram_196__1 (.Q (ram_196__1), .QB (\$dummy [308]), .D (nx38220), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38221 (.Y (nx38220), .A0 (ram_196__1), .A1 (nx65920), .S0 (
             nx64188)) ;
    dffr reg_ram_197__1 (.Q (ram_197__1), .QB (\$dummy [309]), .D (nx38210), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38211 (.Y (nx38210), .A0 (ram_197__1), .A1 (nx65920), .S0 (
             nx64184)) ;
    aoi22 ix55850 (.Y (nx55849), .A0 (ram_199__1), .A1 (nx64720), .B0 (
          ram_198__1), .B1 (nx64758)) ;
    dffr reg_ram_199__1 (.Q (ram_199__1), .QB (\$dummy [310]), .D (nx38190), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38191 (.Y (nx38190), .A0 (ram_199__1), .A1 (nx65920), .S0 (
             nx64176)) ;
    dffr reg_ram_198__1 (.Q (ram_198__1), .QB (\$dummy [311]), .D (nx38200), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38201 (.Y (nx38200), .A0 (ram_198__1), .A1 (nx65920), .S0 (
             nx64180)) ;
    nand04 ix6839 (.Y (nx6838), .A0 (nx55858), .A1 (nx55866), .A2 (nx55874), .A3 (
           nx55882)) ;
    aoi22 ix55859 (.Y (nx55858), .A0 (ram_200__1), .A1 (nx64796), .B0 (
          ram_201__1), .B1 (nx64834)) ;
    dffr reg_ram_200__1 (.Q (ram_200__1), .QB (\$dummy [312]), .D (nx38180), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38181 (.Y (nx38180), .A0 (ram_200__1), .A1 (nx65922), .S0 (
             nx64172)) ;
    dffr reg_ram_201__1 (.Q (ram_201__1), .QB (\$dummy [313]), .D (nx38170), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38171 (.Y (nx38170), .A0 (ram_201__1), .A1 (nx65922), .S0 (
             nx64168)) ;
    aoi22 ix55867 (.Y (nx55866), .A0 (ram_203__1), .A1 (nx64872), .B0 (
          ram_202__1), .B1 (nx64910)) ;
    dffr reg_ram_203__1 (.Q (ram_203__1), .QB (\$dummy [314]), .D (nx38150), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38151 (.Y (nx38150), .A0 (ram_203__1), .A1 (nx65922), .S0 (
             nx64160)) ;
    dffr reg_ram_202__1 (.Q (ram_202__1), .QB (\$dummy [315]), .D (nx38160), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38161 (.Y (nx38160), .A0 (ram_202__1), .A1 (nx65922), .S0 (
             nx64164)) ;
    aoi22 ix55875 (.Y (nx55874), .A0 (ram_204__1), .A1 (nx64948), .B0 (
          ram_205__1), .B1 (nx64986)) ;
    dffr reg_ram_204__1 (.Q (ram_204__1), .QB (\$dummy [316]), .D (nx38140), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38141 (.Y (nx38140), .A0 (ram_204__1), .A1 (nx65922), .S0 (
             nx64156)) ;
    dffr reg_ram_205__1 (.Q (ram_205__1), .QB (\$dummy [317]), .D (nx38130), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38131 (.Y (nx38130), .A0 (ram_205__1), .A1 (nx65922), .S0 (
             nx64152)) ;
    aoi22 ix55883 (.Y (nx55882), .A0 (ram_207__1), .A1 (nx65024), .B0 (
          ram_206__1), .B1 (nx65062)) ;
    dffr reg_ram_207__1 (.Q (ram_207__1), .QB (\$dummy [318]), .D (nx38110), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38111 (.Y (nx38110), .A0 (ram_207__1), .A1 (nx65922), .S0 (
             nx64144)) ;
    dffr reg_ram_206__1 (.Q (ram_206__1), .QB (\$dummy [319]), .D (nx38120), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38121 (.Y (nx38120), .A0 (ram_206__1), .A1 (nx65924), .S0 (
             nx64148)) ;
    nand04 ix6761 (.Y (nx6760), .A0 (nx55891), .A1 (nx55959), .A2 (nx56027), .A3 (
           nx56095)) ;
    oai21 ix55892 (.Y (nx55891), .A0 (nx6750), .A1 (nx6672), .B0 (nx65112)) ;
    nand04 ix6751 (.Y (nx6750), .A0 (nx55894), .A1 (nx55902), .A2 (nx55910), .A3 (
           nx55918)) ;
    aoi22 ix55895 (.Y (nx55894), .A0 (ram_80__1), .A1 (nx64494), .B0 (ram_81__1)
          , .B1 (nx64532)) ;
    dffr reg_ram_80__1 (.Q (ram_80__1), .QB (\$dummy [320]), .D (nx38100), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38101 (.Y (nx38100), .A0 (ram_80__1), .A1 (nx65924), .S0 (nx64134
             )) ;
    dffr reg_ram_81__1 (.Q (ram_81__1), .QB (\$dummy [321]), .D (nx38090), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38091 (.Y (nx38090), .A0 (ram_81__1), .A1 (nx65924), .S0 (nx64130
             )) ;
    aoi22 ix55903 (.Y (nx55902), .A0 (ram_83__1), .A1 (nx64570), .B0 (ram_82__1)
          , .B1 (nx64608)) ;
    dffr reg_ram_83__1 (.Q (ram_83__1), .QB (\$dummy [322]), .D (nx38070), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38071 (.Y (nx38070), .A0 (ram_83__1), .A1 (nx65924), .S0 (nx64122
             )) ;
    dffr reg_ram_82__1 (.Q (ram_82__1), .QB (\$dummy [323]), .D (nx38080), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38081 (.Y (nx38080), .A0 (ram_82__1), .A1 (nx65924), .S0 (nx64126
             )) ;
    aoi22 ix55911 (.Y (nx55910), .A0 (ram_84__1), .A1 (nx64646), .B0 (ram_85__1)
          , .B1 (nx64684)) ;
    dffr reg_ram_84__1 (.Q (ram_84__1), .QB (\$dummy [324]), .D (nx38060), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38061 (.Y (nx38060), .A0 (ram_84__1), .A1 (nx65924), .S0 (nx64118
             )) ;
    dffr reg_ram_85__1 (.Q (ram_85__1), .QB (\$dummy [325]), .D (nx38050), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38051 (.Y (nx38050), .A0 (ram_85__1), .A1 (nx65924), .S0 (nx64114
             )) ;
    aoi22 ix55919 (.Y (nx55918), .A0 (ram_87__1), .A1 (nx64722), .B0 (ram_86__1)
          , .B1 (nx64760)) ;
    dffr reg_ram_87__1 (.Q (ram_87__1), .QB (\$dummy [326]), .D (nx38030), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38031 (.Y (nx38030), .A0 (ram_87__1), .A1 (nx65926), .S0 (nx64106
             )) ;
    dffr reg_ram_86__1 (.Q (ram_86__1), .QB (\$dummy [327]), .D (nx38040), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38041 (.Y (nx38040), .A0 (ram_86__1), .A1 (nx65926), .S0 (nx64110
             )) ;
    nand04 ix6673 (.Y (nx6672), .A0 (nx55927), .A1 (nx55935), .A2 (nx55943), .A3 (
           nx55951)) ;
    aoi22 ix55928 (.Y (nx55927), .A0 (ram_88__1), .A1 (nx64798), .B0 (ram_89__1)
          , .B1 (nx64836)) ;
    dffr reg_ram_88__1 (.Q (ram_88__1), .QB (\$dummy [328]), .D (nx38020), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38021 (.Y (nx38020), .A0 (ram_88__1), .A1 (nx65926), .S0 (nx64102
             )) ;
    dffr reg_ram_89__1 (.Q (ram_89__1), .QB (\$dummy [329]), .D (nx38010), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38011 (.Y (nx38010), .A0 (ram_89__1), .A1 (nx65926), .S0 (nx64098
             )) ;
    aoi22 ix55936 (.Y (nx55935), .A0 (ram_91__1), .A1 (nx64874), .B0 (ram_90__1)
          , .B1 (nx64912)) ;
    dffr reg_ram_91__1 (.Q (ram_91__1), .QB (\$dummy [330]), .D (nx37990), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37991 (.Y (nx37990), .A0 (ram_91__1), .A1 (nx65926), .S0 (nx64090
             )) ;
    dffr reg_ram_90__1 (.Q (ram_90__1), .QB (\$dummy [331]), .D (nx38000), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38001 (.Y (nx38000), .A0 (ram_90__1), .A1 (nx65926), .S0 (nx64094
             )) ;
    aoi22 ix55944 (.Y (nx55943), .A0 (ram_92__1), .A1 (nx64950), .B0 (ram_93__1)
          , .B1 (nx64988)) ;
    dffr reg_ram_92__1 (.Q (ram_92__1), .QB (\$dummy [332]), .D (nx37980), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37981 (.Y (nx37980), .A0 (ram_92__1), .A1 (nx65926), .S0 (nx64086
             )) ;
    dffr reg_ram_93__1 (.Q (ram_93__1), .QB (\$dummy [333]), .D (nx37970), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37971 (.Y (nx37970), .A0 (ram_93__1), .A1 (nx65928), .S0 (nx64082
             )) ;
    aoi22 ix55952 (.Y (nx55951), .A0 (ram_95__1), .A1 (nx65026), .B0 (ram_94__1)
          , .B1 (nx65064)) ;
    dffr reg_ram_95__1 (.Q (ram_95__1), .QB (\$dummy [334]), .D (nx37950), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37951 (.Y (nx37950), .A0 (ram_95__1), .A1 (nx65928), .S0 (nx64074
             )) ;
    dffr reg_ram_94__1 (.Q (ram_94__1), .QB (\$dummy [335]), .D (nx37960), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37961 (.Y (nx37960), .A0 (ram_94__1), .A1 (nx65928), .S0 (nx64078
             )) ;
    oai21 ix55960 (.Y (nx55959), .A0 (nx6588), .A1 (nx6510), .B0 (nx65116)) ;
    nand04 ix6589 (.Y (nx6588), .A0 (nx55962), .A1 (nx55970), .A2 (nx55978), .A3 (
           nx55986)) ;
    aoi22 ix55963 (.Y (nx55962), .A0 (ram_64__1), .A1 (nx64494), .B0 (ram_65__1)
          , .B1 (nx64532)) ;
    dffr reg_ram_64__1 (.Q (ram_64__1), .QB (\$dummy [336]), .D (nx37940), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37941 (.Y (nx37940), .A0 (ram_64__1), .A1 (nx65928), .S0 (nx64064
             )) ;
    dffr reg_ram_65__1 (.Q (ram_65__1), .QB (\$dummy [337]), .D (nx37930), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37931 (.Y (nx37930), .A0 (ram_65__1), .A1 (nx65928), .S0 (nx64060
             )) ;
    aoi22 ix55971 (.Y (nx55970), .A0 (ram_67__1), .A1 (nx64570), .B0 (ram_66__1)
          , .B1 (nx64608)) ;
    dffr reg_ram_67__1 (.Q (ram_67__1), .QB (\$dummy [338]), .D (nx37910), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37911 (.Y (nx37910), .A0 (ram_67__1), .A1 (nx65928), .S0 (nx64052
             )) ;
    dffr reg_ram_66__1 (.Q (ram_66__1), .QB (\$dummy [339]), .D (nx37920), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37921 (.Y (nx37920), .A0 (ram_66__1), .A1 (nx65928), .S0 (nx64056
             )) ;
    aoi22 ix55979 (.Y (nx55978), .A0 (ram_68__1), .A1 (nx64646), .B0 (ram_69__1)
          , .B1 (nx64684)) ;
    dffr reg_ram_68__1 (.Q (ram_68__1), .QB (\$dummy [340]), .D (nx37900), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37901 (.Y (nx37900), .A0 (ram_68__1), .A1 (nx65930), .S0 (nx64048
             )) ;
    dffr reg_ram_69__1 (.Q (ram_69__1), .QB (\$dummy [341]), .D (nx37890), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37891 (.Y (nx37890), .A0 (ram_69__1), .A1 (nx65930), .S0 (nx64044
             )) ;
    aoi22 ix55987 (.Y (nx55986), .A0 (ram_71__1), .A1 (nx64722), .B0 (ram_70__1)
          , .B1 (nx64760)) ;
    dffr reg_ram_71__1 (.Q (ram_71__1), .QB (\$dummy [342]), .D (nx37870), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37871 (.Y (nx37870), .A0 (ram_71__1), .A1 (nx65930), .S0 (nx64036
             )) ;
    dffr reg_ram_70__1 (.Q (ram_70__1), .QB (\$dummy [343]), .D (nx37880), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37881 (.Y (nx37880), .A0 (ram_70__1), .A1 (nx65930), .S0 (nx64040
             )) ;
    nand04 ix6511 (.Y (nx6510), .A0 (nx55995), .A1 (nx56003), .A2 (nx56011), .A3 (
           nx56019)) ;
    aoi22 ix55996 (.Y (nx55995), .A0 (ram_72__1), .A1 (nx64798), .B0 (ram_73__1)
          , .B1 (nx64836)) ;
    dffr reg_ram_72__1 (.Q (ram_72__1), .QB (\$dummy [344]), .D (nx37860), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37861 (.Y (nx37860), .A0 (ram_72__1), .A1 (nx65930), .S0 (nx64032
             )) ;
    dffr reg_ram_73__1 (.Q (ram_73__1), .QB (\$dummy [345]), .D (nx37850), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37851 (.Y (nx37850), .A0 (ram_73__1), .A1 (nx65930), .S0 (nx64028
             )) ;
    aoi22 ix56004 (.Y (nx56003), .A0 (ram_75__1), .A1 (nx64874), .B0 (ram_74__1)
          , .B1 (nx64912)) ;
    dffr reg_ram_75__1 (.Q (ram_75__1), .QB (\$dummy [346]), .D (nx37830), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37831 (.Y (nx37830), .A0 (ram_75__1), .A1 (nx65930), .S0 (nx64020
             )) ;
    dffr reg_ram_74__1 (.Q (ram_74__1), .QB (\$dummy [347]), .D (nx37840), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37841 (.Y (nx37840), .A0 (ram_74__1), .A1 (nx65932), .S0 (nx64024
             )) ;
    aoi22 ix56012 (.Y (nx56011), .A0 (ram_76__1), .A1 (nx64950), .B0 (ram_77__1)
          , .B1 (nx64988)) ;
    dffr reg_ram_76__1 (.Q (ram_76__1), .QB (\$dummy [348]), .D (nx37820), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37821 (.Y (nx37820), .A0 (ram_76__1), .A1 (nx65932), .S0 (nx64016
             )) ;
    dffr reg_ram_77__1 (.Q (ram_77__1), .QB (\$dummy [349]), .D (nx37810), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37811 (.Y (nx37810), .A0 (ram_77__1), .A1 (nx65932), .S0 (nx64012
             )) ;
    aoi22 ix56020 (.Y (nx56019), .A0 (ram_79__1), .A1 (nx65026), .B0 (ram_78__1)
          , .B1 (nx65064)) ;
    dffr reg_ram_79__1 (.Q (ram_79__1), .QB (\$dummy [350]), .D (nx37790), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37791 (.Y (nx37790), .A0 (ram_79__1), .A1 (nx65932), .S0 (nx64004
             )) ;
    dffr reg_ram_78__1 (.Q (ram_78__1), .QB (\$dummy [351]), .D (nx37800), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37801 (.Y (nx37800), .A0 (ram_78__1), .A1 (nx65932), .S0 (nx64008
             )) ;
    oai21 ix56028 (.Y (nx56027), .A0 (nx6424), .A1 (nx6346), .B0 (nx65120)) ;
    nand04 ix6425 (.Y (nx6424), .A0 (nx56030), .A1 (nx56038), .A2 (nx56046), .A3 (
           nx56054)) ;
    aoi22 ix56031 (.Y (nx56030), .A0 (ram_48__1), .A1 (nx64494), .B0 (ram_49__1)
          , .B1 (nx64532)) ;
    dffr reg_ram_48__1 (.Q (ram_48__1), .QB (\$dummy [352]), .D (nx37780), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37781 (.Y (nx37780), .A0 (ram_48__1), .A1 (nx65932), .S0 (nx63994
             )) ;
    dffr reg_ram_49__1 (.Q (ram_49__1), .QB (\$dummy [353]), .D (nx37770), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37771 (.Y (nx37770), .A0 (ram_49__1), .A1 (nx65932), .S0 (nx63990
             )) ;
    aoi22 ix56039 (.Y (nx56038), .A0 (ram_51__1), .A1 (nx64570), .B0 (ram_50__1)
          , .B1 (nx64608)) ;
    dffr reg_ram_51__1 (.Q (ram_51__1), .QB (\$dummy [354]), .D (nx37750), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37751 (.Y (nx37750), .A0 (ram_51__1), .A1 (nx65934), .S0 (nx63982
             )) ;
    dffr reg_ram_50__1 (.Q (ram_50__1), .QB (\$dummy [355]), .D (nx37760), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37761 (.Y (nx37760), .A0 (ram_50__1), .A1 (nx65934), .S0 (nx63986
             )) ;
    aoi22 ix56047 (.Y (nx56046), .A0 (ram_52__1), .A1 (nx64646), .B0 (ram_53__1)
          , .B1 (nx64684)) ;
    dffr reg_ram_52__1 (.Q (ram_52__1), .QB (\$dummy [356]), .D (nx37740), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37741 (.Y (nx37740), .A0 (ram_52__1), .A1 (nx65934), .S0 (nx63978
             )) ;
    dffr reg_ram_53__1 (.Q (ram_53__1), .QB (\$dummy [357]), .D (nx37730), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37731 (.Y (nx37730), .A0 (ram_53__1), .A1 (nx65934), .S0 (nx63974
             )) ;
    aoi22 ix56055 (.Y (nx56054), .A0 (ram_55__1), .A1 (nx64722), .B0 (ram_54__1)
          , .B1 (nx64760)) ;
    dffr reg_ram_55__1 (.Q (ram_55__1), .QB (\$dummy [358]), .D (nx37710), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37711 (.Y (nx37710), .A0 (ram_55__1), .A1 (nx65934), .S0 (nx63966
             )) ;
    dffr reg_ram_54__1 (.Q (ram_54__1), .QB (\$dummy [359]), .D (nx37720), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37721 (.Y (nx37720), .A0 (ram_54__1), .A1 (nx65934), .S0 (nx63970
             )) ;
    nand04 ix6347 (.Y (nx6346), .A0 (nx56063), .A1 (nx56071), .A2 (nx56079), .A3 (
           nx56087)) ;
    aoi22 ix56064 (.Y (nx56063), .A0 (ram_56__1), .A1 (nx64798), .B0 (ram_57__1)
          , .B1 (nx64836)) ;
    dffr reg_ram_56__1 (.Q (ram_56__1), .QB (\$dummy [360]), .D (nx37700), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37701 (.Y (nx37700), .A0 (ram_56__1), .A1 (nx65934), .S0 (nx63962
             )) ;
    dffr reg_ram_57__1 (.Q (ram_57__1), .QB (\$dummy [361]), .D (nx37690), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37691 (.Y (nx37690), .A0 (ram_57__1), .A1 (nx65936), .S0 (nx63958
             )) ;
    aoi22 ix56072 (.Y (nx56071), .A0 (ram_59__1), .A1 (nx64874), .B0 (ram_58__1)
          , .B1 (nx64912)) ;
    dffr reg_ram_59__1 (.Q (ram_59__1), .QB (\$dummy [362]), .D (nx37670), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37671 (.Y (nx37670), .A0 (ram_59__1), .A1 (nx65936), .S0 (nx63950
             )) ;
    dffr reg_ram_58__1 (.Q (ram_58__1), .QB (\$dummy [363]), .D (nx37680), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37681 (.Y (nx37680), .A0 (ram_58__1), .A1 (nx65936), .S0 (nx63954
             )) ;
    aoi22 ix56080 (.Y (nx56079), .A0 (ram_60__1), .A1 (nx64950), .B0 (ram_61__1)
          , .B1 (nx64988)) ;
    dffr reg_ram_60__1 (.Q (ram_60__1), .QB (\$dummy [364]), .D (nx37660), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37661 (.Y (nx37660), .A0 (ram_60__1), .A1 (nx65936), .S0 (nx63946
             )) ;
    dffr reg_ram_61__1 (.Q (ram_61__1), .QB (\$dummy [365]), .D (nx37650), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37651 (.Y (nx37650), .A0 (ram_61__1), .A1 (nx65936), .S0 (nx63942
             )) ;
    aoi22 ix56088 (.Y (nx56087), .A0 (ram_63__1), .A1 (nx65026), .B0 (ram_62__1)
          , .B1 (nx65064)) ;
    dffr reg_ram_63__1 (.Q (ram_63__1), .QB (\$dummy [366]), .D (nx37630), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37631 (.Y (nx37630), .A0 (ram_63__1), .A1 (nx65936), .S0 (nx63934
             )) ;
    dffr reg_ram_62__1 (.Q (ram_62__1), .QB (\$dummy [367]), .D (nx37640), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37641 (.Y (nx37640), .A0 (ram_62__1), .A1 (nx65936), .S0 (nx63938
             )) ;
    oai21 ix56096 (.Y (nx56095), .A0 (nx6262), .A1 (nx6184), .B0 (nx65124)) ;
    nand04 ix6263 (.Y (nx6262), .A0 (nx56098), .A1 (nx56106), .A2 (nx56114), .A3 (
           nx56122)) ;
    aoi22 ix56099 (.Y (nx56098), .A0 (ram_32__1), .A1 (nx64494), .B0 (ram_33__1)
          , .B1 (nx64532)) ;
    dffr reg_ram_32__1 (.Q (ram_32__1), .QB (\$dummy [368]), .D (nx37620), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37621 (.Y (nx37620), .A0 (ram_32__1), .A1 (nx65938), .S0 (nx63924
             )) ;
    dffr reg_ram_33__1 (.Q (ram_33__1), .QB (\$dummy [369]), .D (nx37610), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37611 (.Y (nx37610), .A0 (ram_33__1), .A1 (nx65938), .S0 (nx63920
             )) ;
    aoi22 ix56107 (.Y (nx56106), .A0 (ram_35__1), .A1 (nx64570), .B0 (ram_34__1)
          , .B1 (nx64608)) ;
    dffr reg_ram_35__1 (.Q (ram_35__1), .QB (\$dummy [370]), .D (nx37590), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37591 (.Y (nx37590), .A0 (ram_35__1), .A1 (nx65938), .S0 (nx63912
             )) ;
    dffr reg_ram_34__1 (.Q (ram_34__1), .QB (\$dummy [371]), .D (nx37600), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37601 (.Y (nx37600), .A0 (ram_34__1), .A1 (nx65938), .S0 (nx63916
             )) ;
    aoi22 ix56115 (.Y (nx56114), .A0 (ram_36__1), .A1 (nx64646), .B0 (ram_37__1)
          , .B1 (nx64684)) ;
    dffr reg_ram_36__1 (.Q (ram_36__1), .QB (\$dummy [372]), .D (nx37580), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37581 (.Y (nx37580), .A0 (ram_36__1), .A1 (nx65938), .S0 (nx63908
             )) ;
    dffr reg_ram_37__1 (.Q (ram_37__1), .QB (\$dummy [373]), .D (nx37570), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37571 (.Y (nx37570), .A0 (ram_37__1), .A1 (nx65938), .S0 (nx63904
             )) ;
    aoi22 ix56123 (.Y (nx56122), .A0 (ram_39__1), .A1 (nx64722), .B0 (ram_38__1)
          , .B1 (nx64760)) ;
    dffr reg_ram_39__1 (.Q (ram_39__1), .QB (\$dummy [374]), .D (nx37550), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37551 (.Y (nx37550), .A0 (ram_39__1), .A1 (nx65938), .S0 (nx63896
             )) ;
    dffr reg_ram_38__1 (.Q (ram_38__1), .QB (\$dummy [375]), .D (nx37560), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37561 (.Y (nx37560), .A0 (ram_38__1), .A1 (nx65940), .S0 (nx63900
             )) ;
    nand04 ix6185 (.Y (nx6184), .A0 (nx56131), .A1 (nx56139), .A2 (nx56147), .A3 (
           nx56155)) ;
    aoi22 ix56132 (.Y (nx56131), .A0 (ram_40__1), .A1 (nx64798), .B0 (ram_41__1)
          , .B1 (nx64836)) ;
    dffr reg_ram_40__1 (.Q (ram_40__1), .QB (\$dummy [376]), .D (nx37540), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37541 (.Y (nx37540), .A0 (ram_40__1), .A1 (nx65940), .S0 (nx63892
             )) ;
    dffr reg_ram_41__1 (.Q (ram_41__1), .QB (\$dummy [377]), .D (nx37530), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37531 (.Y (nx37530), .A0 (ram_41__1), .A1 (nx65940), .S0 (nx63888
             )) ;
    aoi22 ix56140 (.Y (nx56139), .A0 (ram_43__1), .A1 (nx64874), .B0 (ram_42__1)
          , .B1 (nx64912)) ;
    dffr reg_ram_43__1 (.Q (ram_43__1), .QB (\$dummy [378]), .D (nx37510), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37511 (.Y (nx37510), .A0 (ram_43__1), .A1 (nx65940), .S0 (nx63880
             )) ;
    dffr reg_ram_42__1 (.Q (ram_42__1), .QB (\$dummy [379]), .D (nx37520), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37521 (.Y (nx37520), .A0 (ram_42__1), .A1 (nx65940), .S0 (nx63884
             )) ;
    aoi22 ix56148 (.Y (nx56147), .A0 (ram_44__1), .A1 (nx64950), .B0 (ram_45__1)
          , .B1 (nx64988)) ;
    dffr reg_ram_44__1 (.Q (ram_44__1), .QB (\$dummy [380]), .D (nx37500), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37501 (.Y (nx37500), .A0 (ram_44__1), .A1 (nx65940), .S0 (nx63876
             )) ;
    dffr reg_ram_45__1 (.Q (ram_45__1), .QB (\$dummy [381]), .D (nx37490), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37491 (.Y (nx37490), .A0 (ram_45__1), .A1 (nx65940), .S0 (nx63872
             )) ;
    aoi22 ix56156 (.Y (nx56155), .A0 (ram_47__1), .A1 (nx65026), .B0 (ram_46__1)
          , .B1 (nx65064)) ;
    dffr reg_ram_47__1 (.Q (ram_47__1), .QB (\$dummy [382]), .D (nx37470), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37471 (.Y (nx37470), .A0 (ram_47__1), .A1 (nx65942), .S0 (nx63864
             )) ;
    dffr reg_ram_46__1 (.Q (ram_46__1), .QB (\$dummy [383]), .D (nx37480), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37481 (.Y (nx37480), .A0 (ram_46__1), .A1 (nx65942), .S0 (nx63868
             )) ;
    nand04 ix6105 (.Y (nx6104), .A0 (nx56164), .A1 (nx56232), .A2 (nx56300), .A3 (
           nx56368)) ;
    oai21 ix56165 (.Y (nx56164), .A0 (nx6094), .A1 (nx6016), .B0 (nx65128)) ;
    nand04 ix6095 (.Y (nx6094), .A0 (nx56167), .A1 (nx56175), .A2 (nx56183), .A3 (
           nx56191)) ;
    aoi22 ix56168 (.Y (nx56167), .A0 (ram_16__1), .A1 (nx64494), .B0 (ram_17__1)
          , .B1 (nx64532)) ;
    dffr reg_ram_16__1 (.Q (ram_16__1), .QB (\$dummy [384]), .D (nx37460), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37461 (.Y (nx37460), .A0 (ram_16__1), .A1 (nx65942), .S0 (nx63854
             )) ;
    dffr reg_ram_17__1 (.Q (ram_17__1), .QB (\$dummy [385]), .D (nx37450), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37451 (.Y (nx37450), .A0 (ram_17__1), .A1 (nx65942), .S0 (nx63850
             )) ;
    aoi22 ix56176 (.Y (nx56175), .A0 (ram_19__1), .A1 (nx64570), .B0 (ram_18__1)
          , .B1 (nx64608)) ;
    dffr reg_ram_19__1 (.Q (ram_19__1), .QB (\$dummy [386]), .D (nx37430), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37431 (.Y (nx37430), .A0 (ram_19__1), .A1 (nx65942), .S0 (nx63842
             )) ;
    dffr reg_ram_18__1 (.Q (ram_18__1), .QB (\$dummy [387]), .D (nx37440), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37441 (.Y (nx37440), .A0 (ram_18__1), .A1 (nx65942), .S0 (nx63846
             )) ;
    aoi22 ix56184 (.Y (nx56183), .A0 (ram_20__1), .A1 (nx64646), .B0 (ram_21__1)
          , .B1 (nx64684)) ;
    dffr reg_ram_20__1 (.Q (ram_20__1), .QB (\$dummy [388]), .D (nx37420), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37421 (.Y (nx37420), .A0 (ram_20__1), .A1 (nx65942), .S0 (nx63838
             )) ;
    dffr reg_ram_21__1 (.Q (ram_21__1), .QB (\$dummy [389]), .D (nx37410), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37411 (.Y (nx37410), .A0 (ram_21__1), .A1 (nx65944), .S0 (nx63834
             )) ;
    aoi22 ix56192 (.Y (nx56191), .A0 (ram_23__1), .A1 (nx64722), .B0 (ram_22__1)
          , .B1 (nx64760)) ;
    dffr reg_ram_23__1 (.Q (ram_23__1), .QB (\$dummy [390]), .D (nx37390), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37391 (.Y (nx37390), .A0 (ram_23__1), .A1 (nx65944), .S0 (nx63826
             )) ;
    dffr reg_ram_22__1 (.Q (ram_22__1), .QB (\$dummy [391]), .D (nx37400), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37401 (.Y (nx37400), .A0 (ram_22__1), .A1 (nx65944), .S0 (nx63830
             )) ;
    nand04 ix6017 (.Y (nx6016), .A0 (nx56200), .A1 (nx56208), .A2 (nx56216), .A3 (
           nx56224)) ;
    aoi22 ix56201 (.Y (nx56200), .A0 (ram_24__1), .A1 (nx64798), .B0 (ram_25__1)
          , .B1 (nx64836)) ;
    dffr reg_ram_24__1 (.Q (ram_24__1), .QB (\$dummy [392]), .D (nx37380), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37381 (.Y (nx37380), .A0 (ram_24__1), .A1 (nx65944), .S0 (nx63822
             )) ;
    dffr reg_ram_25__1 (.Q (ram_25__1), .QB (\$dummy [393]), .D (nx37370), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37371 (.Y (nx37370), .A0 (ram_25__1), .A1 (nx65944), .S0 (nx63818
             )) ;
    aoi22 ix56209 (.Y (nx56208), .A0 (ram_27__1), .A1 (nx64874), .B0 (ram_26__1)
          , .B1 (nx64912)) ;
    dffr reg_ram_27__1 (.Q (ram_27__1), .QB (\$dummy [394]), .D (nx37350), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37351 (.Y (nx37350), .A0 (ram_27__1), .A1 (nx65944), .S0 (nx63810
             )) ;
    dffr reg_ram_26__1 (.Q (ram_26__1), .QB (\$dummy [395]), .D (nx37360), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37361 (.Y (nx37360), .A0 (ram_26__1), .A1 (nx65944), .S0 (nx63814
             )) ;
    aoi22 ix56217 (.Y (nx56216), .A0 (ram_28__1), .A1 (nx64950), .B0 (ram_29__1)
          , .B1 (nx64988)) ;
    dffr reg_ram_28__1 (.Q (ram_28__1), .QB (\$dummy [396]), .D (nx37340), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37341 (.Y (nx37340), .A0 (ram_28__1), .A1 (nx65946), .S0 (nx63806
             )) ;
    dffr reg_ram_29__1 (.Q (ram_29__1), .QB (\$dummy [397]), .D (nx37330), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37331 (.Y (nx37330), .A0 (ram_29__1), .A1 (nx65946), .S0 (nx63802
             )) ;
    aoi22 ix56225 (.Y (nx56224), .A0 (ram_31__1), .A1 (nx65026), .B0 (ram_30__1)
          , .B1 (nx65064)) ;
    dffr reg_ram_31__1 (.Q (ram_31__1), .QB (\$dummy [398]), .D (nx37310), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37311 (.Y (nx37310), .A0 (ram_31__1), .A1 (nx65946), .S0 (nx63794
             )) ;
    dffr reg_ram_30__1 (.Q (ram_30__1), .QB (\$dummy [399]), .D (nx37320), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37321 (.Y (nx37320), .A0 (ram_30__1), .A1 (nx65946), .S0 (nx63798
             )) ;
    oai21 ix56233 (.Y (nx56232), .A0 (nx5932), .A1 (nx5854), .B0 (nx65142)) ;
    nand04 ix5933 (.Y (nx5932), .A0 (nx56235), .A1 (nx56243), .A2 (nx56251), .A3 (
           nx56259)) ;
    aoi22 ix56236 (.Y (nx56235), .A0 (ram_0__1), .A1 (nx64494), .B0 (ram_1__1), 
          .B1 (nx64532)) ;
    dffr reg_ram_0__1 (.Q (ram_0__1), .QB (\$dummy [400]), .D (nx37300), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37301 (.Y (nx37300), .A0 (nx65946), .A1 (ram_0__1), .S0 (nx65132)
             ) ;
    dffr reg_ram_1__1 (.Q (ram_1__1), .QB (\$dummy [401]), .D (nx37290), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37291 (.Y (nx37290), .A0 (nx65946), .A1 (ram_1__1), .S0 (nx65146)
             ) ;
    aoi22 ix56244 (.Y (nx56243), .A0 (ram_3__1), .A1 (nx64570), .B0 (ram_2__1), 
          .B1 (nx64608)) ;
    dffr reg_ram_3__1 (.Q (ram_3__1), .QB (\$dummy [402]), .D (nx37270), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37271 (.Y (nx37270), .A0 (nx65946), .A1 (ram_3__1), .S0 (nx65150)
             ) ;
    dffr reg_ram_2__1 (.Q (ram_2__1), .QB (\$dummy [403]), .D (nx37280), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37281 (.Y (nx37280), .A0 (nx65948), .A1 (ram_2__1), .S0 (nx65154)
             ) ;
    aoi22 ix56252 (.Y (nx56251), .A0 (ram_4__1), .A1 (nx64646), .B0 (ram_5__1), 
          .B1 (nx64684)) ;
    dffr reg_ram_4__1 (.Q (ram_4__1), .QB (\$dummy [404]), .D (nx37260), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37261 (.Y (nx37260), .A0 (nx65948), .A1 (ram_4__1), .S0 (nx65158)
             ) ;
    dffr reg_ram_5__1 (.Q (ram_5__1), .QB (\$dummy [405]), .D (nx37250), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37251 (.Y (nx37250), .A0 (nx65948), .A1 (ram_5__1), .S0 (nx65162)
             ) ;
    aoi22 ix56260 (.Y (nx56259), .A0 (ram_7__1), .A1 (nx64722), .B0 (ram_6__1), 
          .B1 (nx64760)) ;
    dffr reg_ram_7__1 (.Q (ram_7__1), .QB (\$dummy [406]), .D (nx37230), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37231 (.Y (nx37230), .A0 (nx65948), .A1 (ram_7__1), .S0 (nx65166)
             ) ;
    dffr reg_ram_6__1 (.Q (ram_6__1), .QB (\$dummy [407]), .D (nx37240), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37241 (.Y (nx37240), .A0 (nx65948), .A1 (ram_6__1), .S0 (nx65170)
             ) ;
    nand04 ix5855 (.Y (nx5854), .A0 (nx56268), .A1 (nx56276), .A2 (nx56284), .A3 (
           nx56292)) ;
    aoi22 ix56269 (.Y (nx56268), .A0 (ram_8__1), .A1 (nx64798), .B0 (ram_9__1), 
          .B1 (nx64836)) ;
    dffr reg_ram_8__1 (.Q (ram_8__1), .QB (\$dummy [408]), .D (nx37220), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37221 (.Y (nx37220), .A0 (nx65948), .A1 (ram_8__1), .S0 (nx65174)
             ) ;
    dffr reg_ram_9__1 (.Q (ram_9__1), .QB (\$dummy [409]), .D (nx37210), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37211 (.Y (nx37210), .A0 (nx65948), .A1 (ram_9__1), .S0 (nx65178)
             ) ;
    aoi22 ix56277 (.Y (nx56276), .A0 (ram_11__1), .A1 (nx64874), .B0 (ram_10__1)
          , .B1 (nx64912)) ;
    dffr reg_ram_11__1 (.Q (ram_11__1), .QB (\$dummy [410]), .D (nx37190), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37191 (.Y (nx37190), .A0 (nx65950), .A1 (ram_11__1), .S0 (nx65182
             )) ;
    dffr reg_ram_10__1 (.Q (ram_10__1), .QB (\$dummy [411]), .D (nx37200), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37201 (.Y (nx37200), .A0 (nx65950), .A1 (ram_10__1), .S0 (nx65186
             )) ;
    aoi22 ix56285 (.Y (nx56284), .A0 (ram_12__1), .A1 (nx64950), .B0 (ram_13__1)
          , .B1 (nx64988)) ;
    dffr reg_ram_12__1 (.Q (ram_12__1), .QB (\$dummy [412]), .D (nx37180), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37181 (.Y (nx37180), .A0 (nx65950), .A1 (ram_12__1), .S0 (nx65190
             )) ;
    dffr reg_ram_13__1 (.Q (ram_13__1), .QB (\$dummy [413]), .D (nx37170), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37171 (.Y (nx37170), .A0 (nx65950), .A1 (ram_13__1), .S0 (nx65194
             )) ;
    aoi22 ix56293 (.Y (nx56292), .A0 (ram_15__1), .A1 (nx65026), .B0 (ram_14__1)
          , .B1 (nx65064)) ;
    dffr reg_ram_15__1 (.Q (ram_15__1), .QB (\$dummy [414]), .D (nx37150), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37151 (.Y (nx37150), .A0 (nx65950), .A1 (ram_15__1), .S0 (nx65198
             )) ;
    dffr reg_ram_14__1 (.Q (ram_14__1), .QB (\$dummy [415]), .D (nx37160), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37161 (.Y (nx37160), .A0 (nx65950), .A1 (ram_14__1), .S0 (nx65202
             )) ;
    oai21 ix56301 (.Y (nx56300), .A0 (nx5768), .A1 (nx5690), .B0 (nx65206)) ;
    nand04 ix5769 (.Y (nx5768), .A0 (nx56303), .A1 (nx56311), .A2 (nx56319), .A3 (
           nx56327)) ;
    aoi22 ix56304 (.Y (nx56303), .A0 (ram_96__1), .A1 (nx64494), .B0 (ram_97__1)
          , .B1 (nx64532)) ;
    dffr reg_ram_96__1 (.Q (ram_96__1), .QB (\$dummy [416]), .D (nx37140), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37141 (.Y (nx37140), .A0 (ram_96__1), .A1 (nx65950), .S0 (nx63784
             )) ;
    dffr reg_ram_97__1 (.Q (ram_97__1), .QB (\$dummy [417]), .D (nx37130), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37131 (.Y (nx37130), .A0 (ram_97__1), .A1 (nx65952), .S0 (nx63780
             )) ;
    aoi22 ix56312 (.Y (nx56311), .A0 (ram_99__1), .A1 (nx64570), .B0 (ram_98__1)
          , .B1 (nx64608)) ;
    dffr reg_ram_99__1 (.Q (ram_99__1), .QB (\$dummy [418]), .D (nx37110), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37111 (.Y (nx37110), .A0 (ram_99__1), .A1 (nx65952), .S0 (nx63772
             )) ;
    dffr reg_ram_98__1 (.Q (ram_98__1), .QB (\$dummy [419]), .D (nx37120), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37121 (.Y (nx37120), .A0 (ram_98__1), .A1 (nx65952), .S0 (nx63776
             )) ;
    aoi22 ix56320 (.Y (nx56319), .A0 (ram_100__1), .A1 (nx64646), .B0 (
          ram_101__1), .B1 (nx64684)) ;
    dffr reg_ram_100__1 (.Q (ram_100__1), .QB (\$dummy [420]), .D (nx37100), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37101 (.Y (nx37100), .A0 (ram_100__1), .A1 (nx65952), .S0 (
             nx63768)) ;
    dffr reg_ram_101__1 (.Q (ram_101__1), .QB (\$dummy [421]), .D (nx37090), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37091 (.Y (nx37090), .A0 (ram_101__1), .A1 (nx65952), .S0 (
             nx63764)) ;
    aoi22 ix56328 (.Y (nx56327), .A0 (ram_103__1), .A1 (nx64722), .B0 (
          ram_102__1), .B1 (nx64760)) ;
    dffr reg_ram_103__1 (.Q (ram_103__1), .QB (\$dummy [422]), .D (nx37070), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37071 (.Y (nx37070), .A0 (ram_103__1), .A1 (nx65952), .S0 (
             nx63756)) ;
    dffr reg_ram_102__1 (.Q (ram_102__1), .QB (\$dummy [423]), .D (nx37080), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37081 (.Y (nx37080), .A0 (ram_102__1), .A1 (nx65952), .S0 (
             nx63760)) ;
    nand04 ix5691 (.Y (nx5690), .A0 (nx56336), .A1 (nx56344), .A2 (nx56352), .A3 (
           nx56360)) ;
    aoi22 ix56337 (.Y (nx56336), .A0 (ram_104__1), .A1 (nx64798), .B0 (
          ram_105__1), .B1 (nx64836)) ;
    dffr reg_ram_104__1 (.Q (ram_104__1), .QB (\$dummy [424]), .D (nx37060), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37061 (.Y (nx37060), .A0 (ram_104__1), .A1 (nx65954), .S0 (
             nx63752)) ;
    dffr reg_ram_105__1 (.Q (ram_105__1), .QB (\$dummy [425]), .D (nx37050), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37051 (.Y (nx37050), .A0 (ram_105__1), .A1 (nx65954), .S0 (
             nx63748)) ;
    aoi22 ix56345 (.Y (nx56344), .A0 (ram_107__1), .A1 (nx64874), .B0 (
          ram_106__1), .B1 (nx64912)) ;
    dffr reg_ram_107__1 (.Q (ram_107__1), .QB (\$dummy [426]), .D (nx37030), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37031 (.Y (nx37030), .A0 (ram_107__1), .A1 (nx65954), .S0 (
             nx63740)) ;
    dffr reg_ram_106__1 (.Q (ram_106__1), .QB (\$dummy [427]), .D (nx37040), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37041 (.Y (nx37040), .A0 (ram_106__1), .A1 (nx65954), .S0 (
             nx63744)) ;
    aoi22 ix56353 (.Y (nx56352), .A0 (ram_108__1), .A1 (nx64950), .B0 (
          ram_109__1), .B1 (nx64988)) ;
    dffr reg_ram_108__1 (.Q (ram_108__1), .QB (\$dummy [428]), .D (nx37020), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37021 (.Y (nx37020), .A0 (ram_108__1), .A1 (nx65954), .S0 (
             nx63736)) ;
    dffr reg_ram_109__1 (.Q (ram_109__1), .QB (\$dummy [429]), .D (nx37010), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37011 (.Y (nx37010), .A0 (ram_109__1), .A1 (nx65954), .S0 (
             nx63732)) ;
    aoi22 ix56361 (.Y (nx56360), .A0 (ram_111__1), .A1 (nx65026), .B0 (
          ram_110__1), .B1 (nx65064)) ;
    dffr reg_ram_111__1 (.Q (ram_111__1), .QB (\$dummy [430]), .D (nx36990), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36991 (.Y (nx36990), .A0 (ram_111__1), .A1 (nx65954), .S0 (
             nx63724)) ;
    dffr reg_ram_110__1 (.Q (ram_110__1), .QB (\$dummy [431]), .D (nx37000), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix37001 (.Y (nx37000), .A0 (ram_110__1), .A1 (nx65956), .S0 (
             nx63728)) ;
    oai21 ix56369 (.Y (nx56368), .A0 (nx5606), .A1 (nx5528), .B0 (nx65210)) ;
    nand04 ix5607 (.Y (nx5606), .A0 (nx56371), .A1 (nx56379), .A2 (nx56387), .A3 (
           nx56395)) ;
    aoi22 ix56372 (.Y (nx56371), .A0 (ram_112__1), .A1 (nx64496), .B0 (
          ram_113__1), .B1 (nx64534)) ;
    dffr reg_ram_112__1 (.Q (ram_112__1), .QB (\$dummy [432]), .D (nx36980), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36981 (.Y (nx36980), .A0 (ram_112__1), .A1 (nx65956), .S0 (
             nx63714)) ;
    dffr reg_ram_113__1 (.Q (ram_113__1), .QB (\$dummy [433]), .D (nx36970), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36971 (.Y (nx36970), .A0 (ram_113__1), .A1 (nx65956), .S0 (
             nx63710)) ;
    aoi22 ix56380 (.Y (nx56379), .A0 (ram_115__1), .A1 (nx64572), .B0 (
          ram_114__1), .B1 (nx64610)) ;
    dffr reg_ram_115__1 (.Q (ram_115__1), .QB (\$dummy [434]), .D (nx36950), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36951 (.Y (nx36950), .A0 (ram_115__1), .A1 (nx65956), .S0 (
             nx63702)) ;
    dffr reg_ram_114__1 (.Q (ram_114__1), .QB (\$dummy [435]), .D (nx36960), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36961 (.Y (nx36960), .A0 (ram_114__1), .A1 (nx65956), .S0 (
             nx63706)) ;
    aoi22 ix56388 (.Y (nx56387), .A0 (ram_116__1), .A1 (nx64648), .B0 (
          ram_117__1), .B1 (nx64686)) ;
    dffr reg_ram_116__1 (.Q (ram_116__1), .QB (\$dummy [436]), .D (nx36940), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36941 (.Y (nx36940), .A0 (ram_116__1), .A1 (nx65956), .S0 (
             nx63698)) ;
    dffr reg_ram_117__1 (.Q (ram_117__1), .QB (\$dummy [437]), .D (nx36930), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36931 (.Y (nx36930), .A0 (ram_117__1), .A1 (nx65956), .S0 (
             nx63694)) ;
    aoi22 ix56396 (.Y (nx56395), .A0 (ram_119__1), .A1 (nx64724), .B0 (
          ram_118__1), .B1 (nx64762)) ;
    dffr reg_ram_119__1 (.Q (ram_119__1), .QB (\$dummy [438]), .D (nx36910), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36911 (.Y (nx36910), .A0 (ram_119__1), .A1 (nx65958), .S0 (
             nx63686)) ;
    dffr reg_ram_118__1 (.Q (ram_118__1), .QB (\$dummy [439]), .D (nx36920), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36921 (.Y (nx36920), .A0 (ram_118__1), .A1 (nx65958), .S0 (
             nx63690)) ;
    nand04 ix5529 (.Y (nx5528), .A0 (nx56404), .A1 (nx56412), .A2 (nx56420), .A3 (
           nx56428)) ;
    aoi22 ix56405 (.Y (nx56404), .A0 (ram_120__1), .A1 (nx64800), .B0 (
          ram_121__1), .B1 (nx64838)) ;
    dffr reg_ram_120__1 (.Q (ram_120__1), .QB (\$dummy [440]), .D (nx36900), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36901 (.Y (nx36900), .A0 (ram_120__1), .A1 (nx65958), .S0 (
             nx63682)) ;
    dffr reg_ram_121__1 (.Q (ram_121__1), .QB (\$dummy [441]), .D (nx36890), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36891 (.Y (nx36890), .A0 (ram_121__1), .A1 (nx65958), .S0 (
             nx63678)) ;
    aoi22 ix56413 (.Y (nx56412), .A0 (ram_123__1), .A1 (nx64876), .B0 (
          ram_122__1), .B1 (nx64914)) ;
    dffr reg_ram_123__1 (.Q (ram_123__1), .QB (\$dummy [442]), .D (nx36870), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36871 (.Y (nx36870), .A0 (ram_123__1), .A1 (nx65958), .S0 (
             nx63670)) ;
    dffr reg_ram_122__1 (.Q (ram_122__1), .QB (\$dummy [443]), .D (nx36880), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36881 (.Y (nx36880), .A0 (ram_122__1), .A1 (nx65958), .S0 (
             nx63674)) ;
    aoi22 ix56421 (.Y (nx56420), .A0 (ram_124__1), .A1 (nx64952), .B0 (
          ram_125__1), .B1 (nx64990)) ;
    dffr reg_ram_124__1 (.Q (ram_124__1), .QB (\$dummy [444]), .D (nx36860), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36861 (.Y (nx36860), .A0 (ram_124__1), .A1 (nx65958), .S0 (
             nx63666)) ;
    dffr reg_ram_125__1 (.Q (ram_125__1), .QB (\$dummy [445]), .D (nx36850), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36851 (.Y (nx36850), .A0 (ram_125__1), .A1 (nx65960), .S0 (
             nx63662)) ;
    aoi22 ix56429 (.Y (nx56428), .A0 (ram_127__1), .A1 (nx65028), .B0 (
          ram_126__1), .B1 (nx65066)) ;
    dffr reg_ram_127__1 (.Q (ram_127__1), .QB (\$dummy [446]), .D (nx36830), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36831 (.Y (nx36830), .A0 (ram_127__1), .A1 (nx65960), .S0 (
             nx63654)) ;
    dffr reg_ram_126__1 (.Q (ram_126__1), .QB (\$dummy [447]), .D (nx36840), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36841 (.Y (nx36840), .A0 (ram_126__1), .A1 (nx65960), .S0 (
             nx63658)) ;
    nand04 ix5451 (.Y (nx5450), .A0 (nx56437), .A1 (nx56505), .A2 (nx56573), .A3 (
           nx56641)) ;
    oai21 ix56438 (.Y (nx56437), .A0 (nx5440), .A1 (nx5362), .B0 (nx65214)) ;
    nand04 ix5441 (.Y (nx5440), .A0 (nx56440), .A1 (nx56448), .A2 (nx56456), .A3 (
           nx56464)) ;
    aoi22 ix56441 (.Y (nx56440), .A0 (ram_128__1), .A1 (nx64496), .B0 (
          ram_129__1), .B1 (nx64534)) ;
    dffr reg_ram_128__1 (.Q (ram_128__1), .QB (\$dummy [448]), .D (nx36820), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36821 (.Y (nx36820), .A0 (ram_128__1), .A1 (nx65960), .S0 (
             nx63644)) ;
    dffr reg_ram_129__1 (.Q (ram_129__1), .QB (\$dummy [449]), .D (nx36810), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36811 (.Y (nx36810), .A0 (ram_129__1), .A1 (nx65960), .S0 (
             nx63640)) ;
    aoi22 ix56449 (.Y (nx56448), .A0 (ram_131__1), .A1 (nx64572), .B0 (
          ram_130__1), .B1 (nx64610)) ;
    dffr reg_ram_131__1 (.Q (ram_131__1), .QB (\$dummy [450]), .D (nx36790), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36791 (.Y (nx36790), .A0 (ram_131__1), .A1 (nx65960), .S0 (
             nx63632)) ;
    dffr reg_ram_130__1 (.Q (ram_130__1), .QB (\$dummy [451]), .D (nx36800), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36801 (.Y (nx36800), .A0 (ram_130__1), .A1 (nx65960), .S0 (
             nx63636)) ;
    aoi22 ix56457 (.Y (nx56456), .A0 (ram_132__1), .A1 (nx64648), .B0 (
          ram_133__1), .B1 (nx64686)) ;
    dffr reg_ram_132__1 (.Q (ram_132__1), .QB (\$dummy [452]), .D (nx36780), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36781 (.Y (nx36780), .A0 (ram_132__1), .A1 (nx65962), .S0 (
             nx63628)) ;
    dffr reg_ram_133__1 (.Q (ram_133__1), .QB (\$dummy [453]), .D (nx36770), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36771 (.Y (nx36770), .A0 (ram_133__1), .A1 (nx65962), .S0 (
             nx63624)) ;
    aoi22 ix56465 (.Y (nx56464), .A0 (ram_135__1), .A1 (nx64724), .B0 (
          ram_134__1), .B1 (nx64762)) ;
    dffr reg_ram_135__1 (.Q (ram_135__1), .QB (\$dummy [454]), .D (nx36750), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36751 (.Y (nx36750), .A0 (ram_135__1), .A1 (nx65962), .S0 (
             nx63616)) ;
    dffr reg_ram_134__1 (.Q (ram_134__1), .QB (\$dummy [455]), .D (nx36760), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36761 (.Y (nx36760), .A0 (ram_134__1), .A1 (nx65962), .S0 (
             nx63620)) ;
    nand04 ix5363 (.Y (nx5362), .A0 (nx56473), .A1 (nx56481), .A2 (nx56489), .A3 (
           nx56497)) ;
    aoi22 ix56474 (.Y (nx56473), .A0 (ram_136__1), .A1 (nx64800), .B0 (
          ram_137__1), .B1 (nx64838)) ;
    dffr reg_ram_136__1 (.Q (ram_136__1), .QB (\$dummy [456]), .D (nx36740), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36741 (.Y (nx36740), .A0 (ram_136__1), .A1 (nx65962), .S0 (
             nx63612)) ;
    dffr reg_ram_137__1 (.Q (ram_137__1), .QB (\$dummy [457]), .D (nx36730), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36731 (.Y (nx36730), .A0 (ram_137__1), .A1 (nx65962), .S0 (
             nx63608)) ;
    aoi22 ix56482 (.Y (nx56481), .A0 (ram_139__1), .A1 (nx64876), .B0 (
          ram_138__1), .B1 (nx64914)) ;
    dffr reg_ram_139__1 (.Q (ram_139__1), .QB (\$dummy [458]), .D (nx36710), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36711 (.Y (nx36710), .A0 (ram_139__1), .A1 (nx65962), .S0 (
             nx63600)) ;
    dffr reg_ram_138__1 (.Q (ram_138__1), .QB (\$dummy [459]), .D (nx36720), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36721 (.Y (nx36720), .A0 (ram_138__1), .A1 (nx65964), .S0 (
             nx63604)) ;
    aoi22 ix56490 (.Y (nx56489), .A0 (ram_140__1), .A1 (nx64952), .B0 (
          ram_141__1), .B1 (nx64990)) ;
    dffr reg_ram_140__1 (.Q (ram_140__1), .QB (\$dummy [460]), .D (nx36700), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36701 (.Y (nx36700), .A0 (ram_140__1), .A1 (nx65964), .S0 (
             nx63596)) ;
    dffr reg_ram_141__1 (.Q (ram_141__1), .QB (\$dummy [461]), .D (nx36690), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36691 (.Y (nx36690), .A0 (ram_141__1), .A1 (nx65964), .S0 (
             nx63592)) ;
    aoi22 ix56498 (.Y (nx56497), .A0 (ram_143__1), .A1 (nx65028), .B0 (
          ram_142__1), .B1 (nx65066)) ;
    dffr reg_ram_143__1 (.Q (ram_143__1), .QB (\$dummy [462]), .D (nx36670), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36671 (.Y (nx36670), .A0 (ram_143__1), .A1 (nx65964), .S0 (
             nx63584)) ;
    dffr reg_ram_142__1 (.Q (ram_142__1), .QB (\$dummy [463]), .D (nx36680), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36681 (.Y (nx36680), .A0 (ram_142__1), .A1 (nx65964), .S0 (
             nx63588)) ;
    oai21 ix56506 (.Y (nx56505), .A0 (nx5278), .A1 (nx5200), .B0 (nx65218)) ;
    nand04 ix5279 (.Y (nx5278), .A0 (nx56508), .A1 (nx56516), .A2 (nx56524), .A3 (
           nx56532)) ;
    aoi22 ix56509 (.Y (nx56508), .A0 (ram_144__1), .A1 (nx64496), .B0 (
          ram_145__1), .B1 (nx64534)) ;
    dffr reg_ram_144__1 (.Q (ram_144__1), .QB (\$dummy [464]), .D (nx36660), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36661 (.Y (nx36660), .A0 (ram_144__1), .A1 (nx65964), .S0 (
             nx63574)) ;
    dffr reg_ram_145__1 (.Q (ram_145__1), .QB (\$dummy [465]), .D (nx36650), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36651 (.Y (nx36650), .A0 (ram_145__1), .A1 (nx65964), .S0 (
             nx63570)) ;
    aoi22 ix56517 (.Y (nx56516), .A0 (ram_147__1), .A1 (nx64572), .B0 (
          ram_146__1), .B1 (nx64610)) ;
    dffr reg_ram_147__1 (.Q (ram_147__1), .QB (\$dummy [466]), .D (nx36630), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36631 (.Y (nx36630), .A0 (ram_147__1), .A1 (nx65966), .S0 (
             nx63562)) ;
    dffr reg_ram_146__1 (.Q (ram_146__1), .QB (\$dummy [467]), .D (nx36640), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36641 (.Y (nx36640), .A0 (ram_146__1), .A1 (nx65966), .S0 (
             nx63566)) ;
    aoi22 ix56525 (.Y (nx56524), .A0 (ram_148__1), .A1 (nx64648), .B0 (
          ram_149__1), .B1 (nx64686)) ;
    dffr reg_ram_148__1 (.Q (ram_148__1), .QB (\$dummy [468]), .D (nx36620), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36621 (.Y (nx36620), .A0 (ram_148__1), .A1 (nx65966), .S0 (
             nx63558)) ;
    dffr reg_ram_149__1 (.Q (ram_149__1), .QB (\$dummy [469]), .D (nx36610), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36611 (.Y (nx36610), .A0 (ram_149__1), .A1 (nx65966), .S0 (
             nx63554)) ;
    aoi22 ix56533 (.Y (nx56532), .A0 (ram_151__1), .A1 (nx64724), .B0 (
          ram_150__1), .B1 (nx64762)) ;
    dffr reg_ram_151__1 (.Q (ram_151__1), .QB (\$dummy [470]), .D (nx36590), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36591 (.Y (nx36590), .A0 (ram_151__1), .A1 (nx65966), .S0 (
             nx63546)) ;
    dffr reg_ram_150__1 (.Q (ram_150__1), .QB (\$dummy [471]), .D (nx36600), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36601 (.Y (nx36600), .A0 (ram_150__1), .A1 (nx65966), .S0 (
             nx63550)) ;
    nand04 ix5201 (.Y (nx5200), .A0 (nx56541), .A1 (nx56549), .A2 (nx56557), .A3 (
           nx56565)) ;
    aoi22 ix56542 (.Y (nx56541), .A0 (ram_152__1), .A1 (nx64800), .B0 (
          ram_153__1), .B1 (nx64838)) ;
    dffr reg_ram_152__1 (.Q (ram_152__1), .QB (\$dummy [472]), .D (nx36580), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36581 (.Y (nx36580), .A0 (ram_152__1), .A1 (nx65966), .S0 (
             nx63542)) ;
    dffr reg_ram_153__1 (.Q (ram_153__1), .QB (\$dummy [473]), .D (nx36570), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36571 (.Y (nx36570), .A0 (ram_153__1), .A1 (nx65968), .S0 (
             nx63538)) ;
    aoi22 ix56550 (.Y (nx56549), .A0 (ram_155__1), .A1 (nx64876), .B0 (
          ram_154__1), .B1 (nx64914)) ;
    dffr reg_ram_155__1 (.Q (ram_155__1), .QB (\$dummy [474]), .D (nx36550), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36551 (.Y (nx36550), .A0 (ram_155__1), .A1 (nx65968), .S0 (
             nx63530)) ;
    dffr reg_ram_154__1 (.Q (ram_154__1), .QB (\$dummy [475]), .D (nx36560), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36561 (.Y (nx36560), .A0 (ram_154__1), .A1 (nx65968), .S0 (
             nx63534)) ;
    aoi22 ix56558 (.Y (nx56557), .A0 (ram_156__1), .A1 (nx64952), .B0 (
          ram_157__1), .B1 (nx64990)) ;
    dffr reg_ram_156__1 (.Q (ram_156__1), .QB (\$dummy [476]), .D (nx36540), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36541 (.Y (nx36540), .A0 (ram_156__1), .A1 (nx65968), .S0 (
             nx63526)) ;
    dffr reg_ram_157__1 (.Q (ram_157__1), .QB (\$dummy [477]), .D (nx36530), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36531 (.Y (nx36530), .A0 (ram_157__1), .A1 (nx65968), .S0 (
             nx63522)) ;
    aoi22 ix56566 (.Y (nx56565), .A0 (ram_159__1), .A1 (nx65028), .B0 (
          ram_158__1), .B1 (nx65066)) ;
    dffr reg_ram_159__1 (.Q (ram_159__1), .QB (\$dummy [478]), .D (nx36510), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36511 (.Y (nx36510), .A0 (ram_159__1), .A1 (nx65968), .S0 (
             nx63514)) ;
    dffr reg_ram_158__1 (.Q (ram_158__1), .QB (\$dummy [479]), .D (nx36520), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36521 (.Y (nx36520), .A0 (ram_158__1), .A1 (nx65968), .S0 (
             nx63518)) ;
    oai21 ix56574 (.Y (nx56573), .A0 (nx5114), .A1 (nx5036), .B0 (nx65222)) ;
    nand04 ix5115 (.Y (nx5114), .A0 (nx56576), .A1 (nx56584), .A2 (nx56592), .A3 (
           nx56600)) ;
    aoi22 ix56577 (.Y (nx56576), .A0 (ram_160__1), .A1 (nx64496), .B0 (
          ram_161__1), .B1 (nx64534)) ;
    dffr reg_ram_160__1 (.Q (ram_160__1), .QB (\$dummy [480]), .D (nx36500), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36501 (.Y (nx36500), .A0 (ram_160__1), .A1 (nx65970), .S0 (
             nx63504)) ;
    dffr reg_ram_161__1 (.Q (ram_161__1), .QB (\$dummy [481]), .D (nx36490), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36491 (.Y (nx36490), .A0 (ram_161__1), .A1 (nx65970), .S0 (
             nx63500)) ;
    aoi22 ix56585 (.Y (nx56584), .A0 (ram_163__1), .A1 (nx64572), .B0 (
          ram_162__1), .B1 (nx64610)) ;
    dffr reg_ram_163__1 (.Q (ram_163__1), .QB (\$dummy [482]), .D (nx36470), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36471 (.Y (nx36470), .A0 (ram_163__1), .A1 (nx65970), .S0 (
             nx63492)) ;
    dffr reg_ram_162__1 (.Q (ram_162__1), .QB (\$dummy [483]), .D (nx36480), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36481 (.Y (nx36480), .A0 (ram_162__1), .A1 (nx65970), .S0 (
             nx63496)) ;
    aoi22 ix56593 (.Y (nx56592), .A0 (ram_164__1), .A1 (nx64648), .B0 (
          ram_165__1), .B1 (nx64686)) ;
    dffr reg_ram_164__1 (.Q (ram_164__1), .QB (\$dummy [484]), .D (nx36460), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36461 (.Y (nx36460), .A0 (ram_164__1), .A1 (nx65970), .S0 (
             nx63488)) ;
    dffr reg_ram_165__1 (.Q (ram_165__1), .QB (\$dummy [485]), .D (nx36450), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36451 (.Y (nx36450), .A0 (ram_165__1), .A1 (nx65970), .S0 (
             nx63484)) ;
    aoi22 ix56601 (.Y (nx56600), .A0 (ram_167__1), .A1 (nx64724), .B0 (
          ram_166__1), .B1 (nx64762)) ;
    dffr reg_ram_167__1 (.Q (ram_167__1), .QB (\$dummy [486]), .D (nx36430), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36431 (.Y (nx36430), .A0 (ram_167__1), .A1 (nx65970), .S0 (
             nx63476)) ;
    dffr reg_ram_166__1 (.Q (ram_166__1), .QB (\$dummy [487]), .D (nx36440), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36441 (.Y (nx36440), .A0 (ram_166__1), .A1 (nx65972), .S0 (
             nx63480)) ;
    nand04 ix5037 (.Y (nx5036), .A0 (nx56609), .A1 (nx56617), .A2 (nx56625), .A3 (
           nx56633)) ;
    aoi22 ix56610 (.Y (nx56609), .A0 (ram_168__1), .A1 (nx64800), .B0 (
          ram_169__1), .B1 (nx64838)) ;
    dffr reg_ram_168__1 (.Q (ram_168__1), .QB (\$dummy [488]), .D (nx36420), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36421 (.Y (nx36420), .A0 (ram_168__1), .A1 (nx65972), .S0 (
             nx63472)) ;
    dffr reg_ram_169__1 (.Q (ram_169__1), .QB (\$dummy [489]), .D (nx36410), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36411 (.Y (nx36410), .A0 (ram_169__1), .A1 (nx65972), .S0 (
             nx63468)) ;
    aoi22 ix56618 (.Y (nx56617), .A0 (ram_171__1), .A1 (nx64876), .B0 (
          ram_170__1), .B1 (nx64914)) ;
    dffr reg_ram_171__1 (.Q (ram_171__1), .QB (\$dummy [490]), .D (nx36390), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36391 (.Y (nx36390), .A0 (ram_171__1), .A1 (nx65972), .S0 (
             nx63460)) ;
    dffr reg_ram_170__1 (.Q (ram_170__1), .QB (\$dummy [491]), .D (nx36400), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36401 (.Y (nx36400), .A0 (ram_170__1), .A1 (nx65972), .S0 (
             nx63464)) ;
    aoi22 ix56626 (.Y (nx56625), .A0 (ram_172__1), .A1 (nx64952), .B0 (
          ram_173__1), .B1 (nx64990)) ;
    dffr reg_ram_172__1 (.Q (ram_172__1), .QB (\$dummy [492]), .D (nx36380), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36381 (.Y (nx36380), .A0 (ram_172__1), .A1 (nx65972), .S0 (
             nx63456)) ;
    dffr reg_ram_173__1 (.Q (ram_173__1), .QB (\$dummy [493]), .D (nx36370), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36371 (.Y (nx36370), .A0 (ram_173__1), .A1 (nx65972), .S0 (
             nx63452)) ;
    aoi22 ix56634 (.Y (nx56633), .A0 (ram_175__1), .A1 (nx65028), .B0 (
          ram_174__1), .B1 (nx65066)) ;
    dffr reg_ram_175__1 (.Q (ram_175__1), .QB (\$dummy [494]), .D (nx36350), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36351 (.Y (nx36350), .A0 (ram_175__1), .A1 (nx65974), .S0 (
             nx63444)) ;
    dffr reg_ram_174__1 (.Q (ram_174__1), .QB (\$dummy [495]), .D (nx36360), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36361 (.Y (nx36360), .A0 (ram_174__1), .A1 (nx65974), .S0 (
             nx63448)) ;
    oai21 ix56642 (.Y (nx56641), .A0 (nx4952), .A1 (nx4874), .B0 (nx65226)) ;
    nand04 ix4953 (.Y (nx4952), .A0 (nx56644), .A1 (nx56652), .A2 (nx56660), .A3 (
           nx56668)) ;
    aoi22 ix56645 (.Y (nx56644), .A0 (ram_176__1), .A1 (nx64496), .B0 (
          ram_177__1), .B1 (nx64534)) ;
    dffr reg_ram_176__1 (.Q (ram_176__1), .QB (\$dummy [496]), .D (nx36340), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36341 (.Y (nx36340), .A0 (ram_176__1), .A1 (nx65974), .S0 (
             nx63434)) ;
    dffr reg_ram_177__1 (.Q (ram_177__1), .QB (\$dummy [497]), .D (nx36330), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36331 (.Y (nx36330), .A0 (ram_177__1), .A1 (nx65974), .S0 (
             nx63424)) ;
    aoi22 ix56653 (.Y (nx56652), .A0 (ram_179__1), .A1 (nx64572), .B0 (
          ram_178__1), .B1 (nx64610)) ;
    dffr reg_ram_179__1 (.Q (ram_179__1), .QB (\$dummy [498]), .D (nx36310), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36311 (.Y (nx36310), .A0 (ram_179__1), .A1 (nx65974), .S0 (
             nx63404)) ;
    dffr reg_ram_178__1 (.Q (ram_178__1), .QB (\$dummy [499]), .D (nx36320), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36321 (.Y (nx36320), .A0 (ram_178__1), .A1 (nx65974), .S0 (
             nx63414)) ;
    aoi22 ix56661 (.Y (nx56660), .A0 (ram_180__1), .A1 (nx64648), .B0 (
          ram_181__1), .B1 (nx64686)) ;
    dffr reg_ram_180__1 (.Q (ram_180__1), .QB (\$dummy [500]), .D (nx36300), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36301 (.Y (nx36300), .A0 (ram_180__1), .A1 (nx65974), .S0 (
             nx63394)) ;
    dffr reg_ram_181__1 (.Q (ram_181__1), .QB (\$dummy [501]), .D (nx36290), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36291 (.Y (nx36290), .A0 (ram_181__1), .A1 (nx65976), .S0 (
             nx63384)) ;
    aoi22 ix56669 (.Y (nx56668), .A0 (ram_183__1), .A1 (nx64724), .B0 (
          ram_182__1), .B1 (nx64762)) ;
    dffr reg_ram_183__1 (.Q (ram_183__1), .QB (\$dummy [502]), .D (nx36270), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36271 (.Y (nx36270), .A0 (ram_183__1), .A1 (nx65976), .S0 (
             nx63364)) ;
    dffr reg_ram_182__1 (.Q (ram_182__1), .QB (\$dummy [503]), .D (nx36280), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36281 (.Y (nx36280), .A0 (ram_182__1), .A1 (nx65976), .S0 (
             nx63374)) ;
    nand04 ix4875 (.Y (nx4874), .A0 (nx56677), .A1 (nx56685), .A2 (nx56693), .A3 (
           nx56701)) ;
    aoi22 ix56678 (.Y (nx56677), .A0 (ram_184__1), .A1 (nx64800), .B0 (
          ram_185__1), .B1 (nx64838)) ;
    dffr reg_ram_184__1 (.Q (ram_184__1), .QB (\$dummy [504]), .D (nx36260), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36261 (.Y (nx36260), .A0 (ram_184__1), .A1 (nx65976), .S0 (
             nx63354)) ;
    dffr reg_ram_185__1 (.Q (ram_185__1), .QB (\$dummy [505]), .D (nx36250), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36251 (.Y (nx36250), .A0 (ram_185__1), .A1 (nx65976), .S0 (
             nx63344)) ;
    aoi22 ix56686 (.Y (nx56685), .A0 (ram_187__1), .A1 (nx64876), .B0 (
          ram_186__1), .B1 (nx64914)) ;
    dffr reg_ram_187__1 (.Q (ram_187__1), .QB (\$dummy [506]), .D (nx36230), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36231 (.Y (nx36230), .A0 (ram_187__1), .A1 (nx65976), .S0 (
             nx63324)) ;
    dffr reg_ram_186__1 (.Q (ram_186__1), .QB (\$dummy [507]), .D (nx36240), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36241 (.Y (nx36240), .A0 (ram_186__1), .A1 (nx65976), .S0 (
             nx63334)) ;
    aoi22 ix56694 (.Y (nx56693), .A0 (ram_188__1), .A1 (nx64952), .B0 (
          ram_189__1), .B1 (nx64990)) ;
    dffr reg_ram_188__1 (.Q (ram_188__1), .QB (\$dummy [508]), .D (nx36220), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36221 (.Y (nx36220), .A0 (ram_188__1), .A1 (nx65978), .S0 (
             nx63314)) ;
    dffr reg_ram_189__1 (.Q (ram_189__1), .QB (\$dummy [509]), .D (nx36210), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36211 (.Y (nx36210), .A0 (ram_189__1), .A1 (nx65978), .S0 (
             nx63304)) ;
    aoi22 ix56702 (.Y (nx56701), .A0 (ram_191__1), .A1 (nx65028), .B0 (
          ram_190__1), .B1 (nx65066)) ;
    dffr reg_ram_191__1 (.Q (ram_191__1), .QB (\$dummy [510]), .D (nx36190), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36191 (.Y (nx36190), .A0 (ram_191__1), .A1 (nx65978), .S0 (
             nx63284)) ;
    dffr reg_ram_190__1 (.Q (ram_190__1), .QB (\$dummy [511]), .D (nx36200), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix36201 (.Y (nx36200), .A0 (ram_190__1), .A1 (nx65978), .S0 (
             nx63294)) ;
    or04 ix10041 (.Y (dataout[2]), .A0 (nx10036), .A1 (nx9382), .A2 (nx8726), .A3 (
         nx8072)) ;
    nand04 ix10037 (.Y (nx10036), .A0 (nx56711), .A1 (nx56779), .A2 (nx56847), .A3 (
           nx56915)) ;
    oai21 ix56712 (.Y (nx56711), .A0 (nx10026), .A1 (nx9948), .B0 (nx65096)) ;
    nand04 ix10027 (.Y (nx10026), .A0 (nx56714), .A1 (nx56722), .A2 (nx56730), .A3 (
           nx56738)) ;
    aoi22 ix56715 (.Y (nx56714), .A0 (ram_240__2), .A1 (nx64496), .B0 (
          ram_241__2), .B1 (nx64534)) ;
    dffr reg_ram_240__2 (.Q (ram_240__2), .QB (\$dummy [512]), .D (nx41300), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41301 (.Y (nx41300), .A0 (ram_240__2), .A1 (nx65830), .S0 (
             nx64414)) ;
    dffr reg_ram_241__2 (.Q (ram_241__2), .QB (\$dummy [513]), .D (nx41290), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41291 (.Y (nx41290), .A0 (ram_241__2), .A1 (nx65830), .S0 (
             nx64410)) ;
    aoi22 ix56723 (.Y (nx56722), .A0 (ram_243__2), .A1 (nx64572), .B0 (
          ram_242__2), .B1 (nx64610)) ;
    dffr reg_ram_243__2 (.Q (ram_243__2), .QB (\$dummy [514]), .D (nx41270), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41271 (.Y (nx41270), .A0 (ram_243__2), .A1 (nx65830), .S0 (
             nx64402)) ;
    dffr reg_ram_242__2 (.Q (ram_242__2), .QB (\$dummy [515]), .D (nx41280), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41281 (.Y (nx41280), .A0 (ram_242__2), .A1 (nx65830), .S0 (
             nx64406)) ;
    aoi22 ix56731 (.Y (nx56730), .A0 (ram_244__2), .A1 (nx64648), .B0 (
          ram_245__2), .B1 (nx64686)) ;
    dffr reg_ram_244__2 (.Q (ram_244__2), .QB (\$dummy [516]), .D (nx41260), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41261 (.Y (nx41260), .A0 (ram_244__2), .A1 (nx65830), .S0 (
             nx64398)) ;
    dffr reg_ram_245__2 (.Q (ram_245__2), .QB (\$dummy [517]), .D (nx41250), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41251 (.Y (nx41250), .A0 (ram_245__2), .A1 (nx65830), .S0 (
             nx64394)) ;
    aoi22 ix56739 (.Y (nx56738), .A0 (ram_247__2), .A1 (nx64724), .B0 (
          ram_246__2), .B1 (nx64762)) ;
    dffr reg_ram_247__2 (.Q (ram_247__2), .QB (\$dummy [518]), .D (nx41230), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41231 (.Y (nx41230), .A0 (ram_247__2), .A1 (nx65830), .S0 (
             nx64386)) ;
    dffr reg_ram_246__2 (.Q (ram_246__2), .QB (\$dummy [519]), .D (nx41240), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41241 (.Y (nx41240), .A0 (ram_246__2), .A1 (nx65832), .S0 (
             nx64390)) ;
    nand04 ix9949 (.Y (nx9948), .A0 (nx56747), .A1 (nx56755), .A2 (nx56763), .A3 (
           nx56771)) ;
    aoi22 ix56748 (.Y (nx56747), .A0 (ram_248__2), .A1 (nx64800), .B0 (
          ram_249__2), .B1 (nx64838)) ;
    dffr reg_ram_248__2 (.Q (ram_248__2), .QB (\$dummy [520]), .D (nx41220), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41221 (.Y (nx41220), .A0 (ram_248__2), .A1 (nx65832), .S0 (
             nx64382)) ;
    dffr reg_ram_249__2 (.Q (ram_249__2), .QB (\$dummy [521]), .D (nx41210), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41211 (.Y (nx41210), .A0 (ram_249__2), .A1 (nx65832), .S0 (
             nx64378)) ;
    aoi22 ix56756 (.Y (nx56755), .A0 (ram_251__2), .A1 (nx64876), .B0 (
          ram_250__2), .B1 (nx64914)) ;
    dffr reg_ram_251__2 (.Q (ram_251__2), .QB (\$dummy [522]), .D (nx41190), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41191 (.Y (nx41190), .A0 (ram_251__2), .A1 (nx65832), .S0 (
             nx64370)) ;
    dffr reg_ram_250__2 (.Q (ram_250__2), .QB (\$dummy [523]), .D (nx41200), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41201 (.Y (nx41200), .A0 (ram_250__2), .A1 (nx65832), .S0 (
             nx64374)) ;
    aoi22 ix56764 (.Y (nx56763), .A0 (ram_252__2), .A1 (nx64952), .B0 (
          ram_253__2), .B1 (nx64990)) ;
    dffr reg_ram_252__2 (.Q (ram_252__2), .QB (\$dummy [524]), .D (nx41180), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41181 (.Y (nx41180), .A0 (ram_252__2), .A1 (nx65832), .S0 (
             nx64366)) ;
    dffr reg_ram_253__2 (.Q (ram_253__2), .QB (\$dummy [525]), .D (nx41170), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41171 (.Y (nx41170), .A0 (ram_253__2), .A1 (nx65832), .S0 (
             nx64362)) ;
    aoi22 ix56772 (.Y (nx56771), .A0 (ram_255__2), .A1 (nx65028), .B0 (
          ram_254__2), .B1 (nx65066)) ;
    dffr reg_ram_255__2 (.Q (ram_255__2), .QB (\$dummy [526]), .D (nx41150), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41151 (.Y (nx41150), .A0 (ram_255__2), .A1 (nx65834), .S0 (
             nx64354)) ;
    dffr reg_ram_254__2 (.Q (ram_254__2), .QB (\$dummy [527]), .D (nx41160), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41161 (.Y (nx41160), .A0 (ram_254__2), .A1 (nx65834), .S0 (
             nx64358)) ;
    oai21 ix56780 (.Y (nx56779), .A0 (nx9864), .A1 (nx9786), .B0 (nx65100)) ;
    nand04 ix9865 (.Y (nx9864), .A0 (nx56782), .A1 (nx56790), .A2 (nx56798), .A3 (
           nx56806)) ;
    aoi22 ix56783 (.Y (nx56782), .A0 (ram_224__2), .A1 (nx64496), .B0 (
          ram_225__2), .B1 (nx64534)) ;
    dffr reg_ram_224__2 (.Q (ram_224__2), .QB (\$dummy [528]), .D (nx41140), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41141 (.Y (nx41140), .A0 (ram_224__2), .A1 (nx65834), .S0 (
             nx64344)) ;
    dffr reg_ram_225__2 (.Q (ram_225__2), .QB (\$dummy [529]), .D (nx41130), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41131 (.Y (nx41130), .A0 (ram_225__2), .A1 (nx65834), .S0 (
             nx64340)) ;
    aoi22 ix56791 (.Y (nx56790), .A0 (ram_227__2), .A1 (nx64572), .B0 (
          ram_226__2), .B1 (nx64610)) ;
    dffr reg_ram_227__2 (.Q (ram_227__2), .QB (\$dummy [530]), .D (nx41110), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41111 (.Y (nx41110), .A0 (ram_227__2), .A1 (nx65834), .S0 (
             nx64332)) ;
    dffr reg_ram_226__2 (.Q (ram_226__2), .QB (\$dummy [531]), .D (nx41120), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41121 (.Y (nx41120), .A0 (ram_226__2), .A1 (nx65834), .S0 (
             nx64336)) ;
    aoi22 ix56799 (.Y (nx56798), .A0 (ram_228__2), .A1 (nx64648), .B0 (
          ram_229__2), .B1 (nx64686)) ;
    dffr reg_ram_228__2 (.Q (ram_228__2), .QB (\$dummy [532]), .D (nx41100), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41101 (.Y (nx41100), .A0 (ram_228__2), .A1 (nx65834), .S0 (
             nx64328)) ;
    dffr reg_ram_229__2 (.Q (ram_229__2), .QB (\$dummy [533]), .D (nx41090), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41091 (.Y (nx41090), .A0 (ram_229__2), .A1 (nx65836), .S0 (
             nx64324)) ;
    aoi22 ix56807 (.Y (nx56806), .A0 (ram_231__2), .A1 (nx64724), .B0 (
          ram_230__2), .B1 (nx64762)) ;
    dffr reg_ram_231__2 (.Q (ram_231__2), .QB (\$dummy [534]), .D (nx41070), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41071 (.Y (nx41070), .A0 (ram_231__2), .A1 (nx65836), .S0 (
             nx64316)) ;
    dffr reg_ram_230__2 (.Q (ram_230__2), .QB (\$dummy [535]), .D (nx41080), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41081 (.Y (nx41080), .A0 (ram_230__2), .A1 (nx65836), .S0 (
             nx64320)) ;
    nand04 ix9787 (.Y (nx9786), .A0 (nx56815), .A1 (nx56823), .A2 (nx56831), .A3 (
           nx56839)) ;
    aoi22 ix56816 (.Y (nx56815), .A0 (ram_232__2), .A1 (nx64800), .B0 (
          ram_233__2), .B1 (nx64838)) ;
    dffr reg_ram_232__2 (.Q (ram_232__2), .QB (\$dummy [536]), .D (nx41060), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41061 (.Y (nx41060), .A0 (ram_232__2), .A1 (nx65836), .S0 (
             nx64312)) ;
    dffr reg_ram_233__2 (.Q (ram_233__2), .QB (\$dummy [537]), .D (nx41050), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41051 (.Y (nx41050), .A0 (ram_233__2), .A1 (nx65836), .S0 (
             nx64308)) ;
    aoi22 ix56824 (.Y (nx56823), .A0 (ram_235__2), .A1 (nx64876), .B0 (
          ram_234__2), .B1 (nx64914)) ;
    dffr reg_ram_235__2 (.Q (ram_235__2), .QB (\$dummy [538]), .D (nx41030), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41031 (.Y (nx41030), .A0 (ram_235__2), .A1 (nx65836), .S0 (
             nx64300)) ;
    dffr reg_ram_234__2 (.Q (ram_234__2), .QB (\$dummy [539]), .D (nx41040), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41041 (.Y (nx41040), .A0 (ram_234__2), .A1 (nx65836), .S0 (
             nx64304)) ;
    aoi22 ix56832 (.Y (nx56831), .A0 (ram_236__2), .A1 (nx64952), .B0 (
          ram_237__2), .B1 (nx64990)) ;
    dffr reg_ram_236__2 (.Q (ram_236__2), .QB (\$dummy [540]), .D (nx41020), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41021 (.Y (nx41020), .A0 (ram_236__2), .A1 (nx65838), .S0 (
             nx64296)) ;
    dffr reg_ram_237__2 (.Q (ram_237__2), .QB (\$dummy [541]), .D (nx41010), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41011 (.Y (nx41010), .A0 (ram_237__2), .A1 (nx65838), .S0 (
             nx64292)) ;
    aoi22 ix56840 (.Y (nx56839), .A0 (ram_239__2), .A1 (nx65028), .B0 (
          ram_238__2), .B1 (nx65066)) ;
    dffr reg_ram_239__2 (.Q (ram_239__2), .QB (\$dummy [542]), .D (nx40990), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40991 (.Y (nx40990), .A0 (ram_239__2), .A1 (nx65838), .S0 (
             nx64284)) ;
    dffr reg_ram_238__2 (.Q (ram_238__2), .QB (\$dummy [543]), .D (nx41000), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41001 (.Y (nx41000), .A0 (ram_238__2), .A1 (nx65838), .S0 (
             nx64288)) ;
    oai21 ix56848 (.Y (nx56847), .A0 (nx9700), .A1 (nx9622), .B0 (nx65104)) ;
    nand04 ix9701 (.Y (nx9700), .A0 (nx56850), .A1 (nx56858), .A2 (nx56866), .A3 (
           nx56874)) ;
    aoi22 ix56851 (.Y (nx56850), .A0 (ram_208__2), .A1 (nx64498), .B0 (
          ram_209__2), .B1 (nx64536)) ;
    dffr reg_ram_208__2 (.Q (ram_208__2), .QB (\$dummy [544]), .D (nx40980), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40981 (.Y (nx40980), .A0 (ram_208__2), .A1 (nx65838), .S0 (
             nx64274)) ;
    dffr reg_ram_209__2 (.Q (ram_209__2), .QB (\$dummy [545]), .D (nx40970), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40971 (.Y (nx40970), .A0 (ram_209__2), .A1 (nx65838), .S0 (
             nx64270)) ;
    aoi22 ix56859 (.Y (nx56858), .A0 (ram_211__2), .A1 (nx64574), .B0 (
          ram_210__2), .B1 (nx64612)) ;
    dffr reg_ram_211__2 (.Q (ram_211__2), .QB (\$dummy [546]), .D (nx40950), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40951 (.Y (nx40950), .A0 (ram_211__2), .A1 (nx65838), .S0 (
             nx64262)) ;
    dffr reg_ram_210__2 (.Q (ram_210__2), .QB (\$dummy [547]), .D (nx40960), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40961 (.Y (nx40960), .A0 (ram_210__2), .A1 (nx65840), .S0 (
             nx64266)) ;
    aoi22 ix56867 (.Y (nx56866), .A0 (ram_212__2), .A1 (nx64650), .B0 (
          ram_213__2), .B1 (nx64688)) ;
    dffr reg_ram_212__2 (.Q (ram_212__2), .QB (\$dummy [548]), .D (nx40940), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40941 (.Y (nx40940), .A0 (ram_212__2), .A1 (nx65840), .S0 (
             nx64258)) ;
    dffr reg_ram_213__2 (.Q (ram_213__2), .QB (\$dummy [549]), .D (nx40930), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40931 (.Y (nx40930), .A0 (ram_213__2), .A1 (nx65840), .S0 (
             nx64254)) ;
    aoi22 ix56875 (.Y (nx56874), .A0 (ram_215__2), .A1 (nx64726), .B0 (
          ram_214__2), .B1 (nx64764)) ;
    dffr reg_ram_215__2 (.Q (ram_215__2), .QB (\$dummy [550]), .D (nx40910), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40911 (.Y (nx40910), .A0 (ram_215__2), .A1 (nx65840), .S0 (
             nx64246)) ;
    dffr reg_ram_214__2 (.Q (ram_214__2), .QB (\$dummy [551]), .D (nx40920), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40921 (.Y (nx40920), .A0 (ram_214__2), .A1 (nx65840), .S0 (
             nx64250)) ;
    nand04 ix9623 (.Y (nx9622), .A0 (nx56883), .A1 (nx56891), .A2 (nx56899), .A3 (
           nx56907)) ;
    aoi22 ix56884 (.Y (nx56883), .A0 (ram_216__2), .A1 (nx64802), .B0 (
          ram_217__2), .B1 (nx64840)) ;
    dffr reg_ram_216__2 (.Q (ram_216__2), .QB (\$dummy [552]), .D (nx40900), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40901 (.Y (nx40900), .A0 (ram_216__2), .A1 (nx65840), .S0 (
             nx64242)) ;
    dffr reg_ram_217__2 (.Q (ram_217__2), .QB (\$dummy [553]), .D (nx40890), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40891 (.Y (nx40890), .A0 (ram_217__2), .A1 (nx65840), .S0 (
             nx64238)) ;
    aoi22 ix56892 (.Y (nx56891), .A0 (ram_219__2), .A1 (nx64878), .B0 (
          ram_218__2), .B1 (nx64916)) ;
    dffr reg_ram_219__2 (.Q (ram_219__2), .QB (\$dummy [554]), .D (nx40870), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40871 (.Y (nx40870), .A0 (ram_219__2), .A1 (nx65842), .S0 (
             nx64230)) ;
    dffr reg_ram_218__2 (.Q (ram_218__2), .QB (\$dummy [555]), .D (nx40880), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40881 (.Y (nx40880), .A0 (ram_218__2), .A1 (nx65842), .S0 (
             nx64234)) ;
    aoi22 ix56900 (.Y (nx56899), .A0 (ram_220__2), .A1 (nx64954), .B0 (
          ram_221__2), .B1 (nx64992)) ;
    dffr reg_ram_220__2 (.Q (ram_220__2), .QB (\$dummy [556]), .D (nx40860), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40861 (.Y (nx40860), .A0 (ram_220__2), .A1 (nx65842), .S0 (
             nx64226)) ;
    dffr reg_ram_221__2 (.Q (ram_221__2), .QB (\$dummy [557]), .D (nx40850), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40851 (.Y (nx40850), .A0 (ram_221__2), .A1 (nx65842), .S0 (
             nx64222)) ;
    aoi22 ix56908 (.Y (nx56907), .A0 (ram_223__2), .A1 (nx65030), .B0 (
          ram_222__2), .B1 (nx65068)) ;
    dffr reg_ram_223__2 (.Q (ram_223__2), .QB (\$dummy [558]), .D (nx40830), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40831 (.Y (nx40830), .A0 (ram_223__2), .A1 (nx65842), .S0 (
             nx64214)) ;
    dffr reg_ram_222__2 (.Q (ram_222__2), .QB (\$dummy [559]), .D (nx40840), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40841 (.Y (nx40840), .A0 (ram_222__2), .A1 (nx65842), .S0 (
             nx64218)) ;
    oai21 ix56916 (.Y (nx56915), .A0 (nx9538), .A1 (nx9460), .B0 (nx65108)) ;
    nand04 ix9539 (.Y (nx9538), .A0 (nx56918), .A1 (nx56926), .A2 (nx56934), .A3 (
           nx56942)) ;
    aoi22 ix56919 (.Y (nx56918), .A0 (ram_192__2), .A1 (nx64498), .B0 (
          ram_193__2), .B1 (nx64536)) ;
    dffr reg_ram_192__2 (.Q (ram_192__2), .QB (\$dummy [560]), .D (nx40820), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40821 (.Y (nx40820), .A0 (ram_192__2), .A1 (nx65842), .S0 (
             nx64204)) ;
    dffr reg_ram_193__2 (.Q (ram_193__2), .QB (\$dummy [561]), .D (nx40810), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40811 (.Y (nx40810), .A0 (ram_193__2), .A1 (nx65844), .S0 (
             nx64200)) ;
    aoi22 ix56927 (.Y (nx56926), .A0 (ram_195__2), .A1 (nx64574), .B0 (
          ram_194__2), .B1 (nx64612)) ;
    dffr reg_ram_195__2 (.Q (ram_195__2), .QB (\$dummy [562]), .D (nx40790), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40791 (.Y (nx40790), .A0 (ram_195__2), .A1 (nx65844), .S0 (
             nx64192)) ;
    dffr reg_ram_194__2 (.Q (ram_194__2), .QB (\$dummy [563]), .D (nx40800), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40801 (.Y (nx40800), .A0 (ram_194__2), .A1 (nx65844), .S0 (
             nx64196)) ;
    aoi22 ix56935 (.Y (nx56934), .A0 (ram_196__2), .A1 (nx64650), .B0 (
          ram_197__2), .B1 (nx64688)) ;
    dffr reg_ram_196__2 (.Q (ram_196__2), .QB (\$dummy [564]), .D (nx40780), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40781 (.Y (nx40780), .A0 (ram_196__2), .A1 (nx65844), .S0 (
             nx64188)) ;
    dffr reg_ram_197__2 (.Q (ram_197__2), .QB (\$dummy [565]), .D (nx40770), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40771 (.Y (nx40770), .A0 (ram_197__2), .A1 (nx65844), .S0 (
             nx64184)) ;
    aoi22 ix56943 (.Y (nx56942), .A0 (ram_199__2), .A1 (nx64726), .B0 (
          ram_198__2), .B1 (nx64764)) ;
    dffr reg_ram_199__2 (.Q (ram_199__2), .QB (\$dummy [566]), .D (nx40750), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40751 (.Y (nx40750), .A0 (ram_199__2), .A1 (nx65844), .S0 (
             nx64176)) ;
    dffr reg_ram_198__2 (.Q (ram_198__2), .QB (\$dummy [567]), .D (nx40760), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40761 (.Y (nx40760), .A0 (ram_198__2), .A1 (nx65844), .S0 (
             nx64180)) ;
    nand04 ix9461 (.Y (nx9460), .A0 (nx56951), .A1 (nx56959), .A2 (nx56967), .A3 (
           nx56975)) ;
    aoi22 ix56952 (.Y (nx56951), .A0 (ram_200__2), .A1 (nx64802), .B0 (
          ram_201__2), .B1 (nx64840)) ;
    dffr reg_ram_200__2 (.Q (ram_200__2), .QB (\$dummy [568]), .D (nx40740), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40741 (.Y (nx40740), .A0 (ram_200__2), .A1 (nx65846), .S0 (
             nx64172)) ;
    dffr reg_ram_201__2 (.Q (ram_201__2), .QB (\$dummy [569]), .D (nx40730), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40731 (.Y (nx40730), .A0 (ram_201__2), .A1 (nx65846), .S0 (
             nx64168)) ;
    aoi22 ix56960 (.Y (nx56959), .A0 (ram_203__2), .A1 (nx64878), .B0 (
          ram_202__2), .B1 (nx64916)) ;
    dffr reg_ram_203__2 (.Q (ram_203__2), .QB (\$dummy [570]), .D (nx40710), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40711 (.Y (nx40710), .A0 (ram_203__2), .A1 (nx65846), .S0 (
             nx64160)) ;
    dffr reg_ram_202__2 (.Q (ram_202__2), .QB (\$dummy [571]), .D (nx40720), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40721 (.Y (nx40720), .A0 (ram_202__2), .A1 (nx65846), .S0 (
             nx64164)) ;
    aoi22 ix56968 (.Y (nx56967), .A0 (ram_204__2), .A1 (nx64954), .B0 (
          ram_205__2), .B1 (nx64992)) ;
    dffr reg_ram_204__2 (.Q (ram_204__2), .QB (\$dummy [572]), .D (nx40700), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40701 (.Y (nx40700), .A0 (ram_204__2), .A1 (nx65846), .S0 (
             nx64156)) ;
    dffr reg_ram_205__2 (.Q (ram_205__2), .QB (\$dummy [573]), .D (nx40690), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40691 (.Y (nx40690), .A0 (ram_205__2), .A1 (nx65846), .S0 (
             nx64152)) ;
    aoi22 ix56976 (.Y (nx56975), .A0 (ram_207__2), .A1 (nx65030), .B0 (
          ram_206__2), .B1 (nx65068)) ;
    dffr reg_ram_207__2 (.Q (ram_207__2), .QB (\$dummy [574]), .D (nx40670), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40671 (.Y (nx40670), .A0 (ram_207__2), .A1 (nx65846), .S0 (
             nx64144)) ;
    dffr reg_ram_206__2 (.Q (ram_206__2), .QB (\$dummy [575]), .D (nx40680), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40681 (.Y (nx40680), .A0 (ram_206__2), .A1 (nx65848), .S0 (
             nx64148)) ;
    nand04 ix9383 (.Y (nx9382), .A0 (nx56984), .A1 (nx57052), .A2 (nx57120), .A3 (
           nx57188)) ;
    oai21 ix56985 (.Y (nx56984), .A0 (nx9372), .A1 (nx9294), .B0 (nx65112)) ;
    nand04 ix9373 (.Y (nx9372), .A0 (nx56987), .A1 (nx56995), .A2 (nx57003), .A3 (
           nx57011)) ;
    aoi22 ix56988 (.Y (nx56987), .A0 (ram_80__2), .A1 (nx64498), .B0 (ram_81__2)
          , .B1 (nx64536)) ;
    dffr reg_ram_80__2 (.Q (ram_80__2), .QB (\$dummy [576]), .D (nx40660), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40661 (.Y (nx40660), .A0 (ram_80__2), .A1 (nx65848), .S0 (nx64134
             )) ;
    dffr reg_ram_81__2 (.Q (ram_81__2), .QB (\$dummy [577]), .D (nx40650), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40651 (.Y (nx40650), .A0 (ram_81__2), .A1 (nx65848), .S0 (nx64130
             )) ;
    aoi22 ix56996 (.Y (nx56995), .A0 (ram_83__2), .A1 (nx64574), .B0 (ram_82__2)
          , .B1 (nx64612)) ;
    dffr reg_ram_83__2 (.Q (ram_83__2), .QB (\$dummy [578]), .D (nx40630), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40631 (.Y (nx40630), .A0 (ram_83__2), .A1 (nx65848), .S0 (nx64122
             )) ;
    dffr reg_ram_82__2 (.Q (ram_82__2), .QB (\$dummy [579]), .D (nx40640), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40641 (.Y (nx40640), .A0 (ram_82__2), .A1 (nx65848), .S0 (nx64126
             )) ;
    aoi22 ix57004 (.Y (nx57003), .A0 (ram_84__2), .A1 (nx64650), .B0 (ram_85__2)
          , .B1 (nx64688)) ;
    dffr reg_ram_84__2 (.Q (ram_84__2), .QB (\$dummy [580]), .D (nx40620), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40621 (.Y (nx40620), .A0 (ram_84__2), .A1 (nx65848), .S0 (nx64118
             )) ;
    dffr reg_ram_85__2 (.Q (ram_85__2), .QB (\$dummy [581]), .D (nx40610), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40611 (.Y (nx40610), .A0 (ram_85__2), .A1 (nx65848), .S0 (nx64114
             )) ;
    aoi22 ix57012 (.Y (nx57011), .A0 (ram_87__2), .A1 (nx64726), .B0 (ram_86__2)
          , .B1 (nx64764)) ;
    dffr reg_ram_87__2 (.Q (ram_87__2), .QB (\$dummy [582]), .D (nx40590), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40591 (.Y (nx40590), .A0 (ram_87__2), .A1 (nx65850), .S0 (nx64106
             )) ;
    dffr reg_ram_86__2 (.Q (ram_86__2), .QB (\$dummy [583]), .D (nx40600), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40601 (.Y (nx40600), .A0 (ram_86__2), .A1 (nx65850), .S0 (nx64110
             )) ;
    nand04 ix9295 (.Y (nx9294), .A0 (nx57020), .A1 (nx57028), .A2 (nx57036), .A3 (
           nx57044)) ;
    aoi22 ix57021 (.Y (nx57020), .A0 (ram_88__2), .A1 (nx64802), .B0 (ram_89__2)
          , .B1 (nx64840)) ;
    dffr reg_ram_88__2 (.Q (ram_88__2), .QB (\$dummy [584]), .D (nx40580), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40581 (.Y (nx40580), .A0 (ram_88__2), .A1 (nx65850), .S0 (nx64102
             )) ;
    dffr reg_ram_89__2 (.Q (ram_89__2), .QB (\$dummy [585]), .D (nx40570), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40571 (.Y (nx40570), .A0 (ram_89__2), .A1 (nx65850), .S0 (nx64098
             )) ;
    aoi22 ix57029 (.Y (nx57028), .A0 (ram_91__2), .A1 (nx64878), .B0 (ram_90__2)
          , .B1 (nx64916)) ;
    dffr reg_ram_91__2 (.Q (ram_91__2), .QB (\$dummy [586]), .D (nx40550), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40551 (.Y (nx40550), .A0 (ram_91__2), .A1 (nx65850), .S0 (nx64090
             )) ;
    dffr reg_ram_90__2 (.Q (ram_90__2), .QB (\$dummy [587]), .D (nx40560), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40561 (.Y (nx40560), .A0 (ram_90__2), .A1 (nx65850), .S0 (nx64094
             )) ;
    aoi22 ix57037 (.Y (nx57036), .A0 (ram_92__2), .A1 (nx64954), .B0 (ram_93__2)
          , .B1 (nx64992)) ;
    dffr reg_ram_92__2 (.Q (ram_92__2), .QB (\$dummy [588]), .D (nx40540), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40541 (.Y (nx40540), .A0 (ram_92__2), .A1 (nx65850), .S0 (nx64086
             )) ;
    dffr reg_ram_93__2 (.Q (ram_93__2), .QB (\$dummy [589]), .D (nx40530), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40531 (.Y (nx40530), .A0 (ram_93__2), .A1 (nx65852), .S0 (nx64082
             )) ;
    aoi22 ix57045 (.Y (nx57044), .A0 (ram_95__2), .A1 (nx65030), .B0 (ram_94__2)
          , .B1 (nx65068)) ;
    dffr reg_ram_95__2 (.Q (ram_95__2), .QB (\$dummy [590]), .D (nx40510), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40511 (.Y (nx40510), .A0 (ram_95__2), .A1 (nx65852), .S0 (nx64074
             )) ;
    dffr reg_ram_94__2 (.Q (ram_94__2), .QB (\$dummy [591]), .D (nx40520), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40521 (.Y (nx40520), .A0 (ram_94__2), .A1 (nx65852), .S0 (nx64078
             )) ;
    oai21 ix57053 (.Y (nx57052), .A0 (nx9210), .A1 (nx9132), .B0 (nx65116)) ;
    nand04 ix9211 (.Y (nx9210), .A0 (nx57055), .A1 (nx57063), .A2 (nx57071), .A3 (
           nx57079)) ;
    aoi22 ix57056 (.Y (nx57055), .A0 (ram_64__2), .A1 (nx64498), .B0 (ram_65__2)
          , .B1 (nx64536)) ;
    dffr reg_ram_64__2 (.Q (ram_64__2), .QB (\$dummy [592]), .D (nx40500), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40501 (.Y (nx40500), .A0 (ram_64__2), .A1 (nx65852), .S0 (nx64064
             )) ;
    dffr reg_ram_65__2 (.Q (ram_65__2), .QB (\$dummy [593]), .D (nx40490), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40491 (.Y (nx40490), .A0 (ram_65__2), .A1 (nx65852), .S0 (nx64060
             )) ;
    aoi22 ix57064 (.Y (nx57063), .A0 (ram_67__2), .A1 (nx64574), .B0 (ram_66__2)
          , .B1 (nx64612)) ;
    dffr reg_ram_67__2 (.Q (ram_67__2), .QB (\$dummy [594]), .D (nx40470), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40471 (.Y (nx40470), .A0 (ram_67__2), .A1 (nx65852), .S0 (nx64052
             )) ;
    dffr reg_ram_66__2 (.Q (ram_66__2), .QB (\$dummy [595]), .D (nx40480), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40481 (.Y (nx40480), .A0 (ram_66__2), .A1 (nx65852), .S0 (nx64056
             )) ;
    aoi22 ix57072 (.Y (nx57071), .A0 (ram_68__2), .A1 (nx64650), .B0 (ram_69__2)
          , .B1 (nx64688)) ;
    dffr reg_ram_68__2 (.Q (ram_68__2), .QB (\$dummy [596]), .D (nx40460), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40461 (.Y (nx40460), .A0 (ram_68__2), .A1 (nx65854), .S0 (nx64048
             )) ;
    dffr reg_ram_69__2 (.Q (ram_69__2), .QB (\$dummy [597]), .D (nx40450), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40451 (.Y (nx40450), .A0 (ram_69__2), .A1 (nx65854), .S0 (nx64044
             )) ;
    aoi22 ix57080 (.Y (nx57079), .A0 (ram_71__2), .A1 (nx64726), .B0 (ram_70__2)
          , .B1 (nx64764)) ;
    dffr reg_ram_71__2 (.Q (ram_71__2), .QB (\$dummy [598]), .D (nx40430), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40431 (.Y (nx40430), .A0 (ram_71__2), .A1 (nx65854), .S0 (nx64036
             )) ;
    dffr reg_ram_70__2 (.Q (ram_70__2), .QB (\$dummy [599]), .D (nx40440), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40441 (.Y (nx40440), .A0 (ram_70__2), .A1 (nx65854), .S0 (nx64040
             )) ;
    nand04 ix9133 (.Y (nx9132), .A0 (nx57088), .A1 (nx57096), .A2 (nx57104), .A3 (
           nx57112)) ;
    aoi22 ix57089 (.Y (nx57088), .A0 (ram_72__2), .A1 (nx64802), .B0 (ram_73__2)
          , .B1 (nx64840)) ;
    dffr reg_ram_72__2 (.Q (ram_72__2), .QB (\$dummy [600]), .D (nx40420), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40421 (.Y (nx40420), .A0 (ram_72__2), .A1 (nx65854), .S0 (nx64032
             )) ;
    dffr reg_ram_73__2 (.Q (ram_73__2), .QB (\$dummy [601]), .D (nx40410), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40411 (.Y (nx40410), .A0 (ram_73__2), .A1 (nx65854), .S0 (nx64028
             )) ;
    aoi22 ix57097 (.Y (nx57096), .A0 (ram_75__2), .A1 (nx64878), .B0 (ram_74__2)
          , .B1 (nx64916)) ;
    dffr reg_ram_75__2 (.Q (ram_75__2), .QB (\$dummy [602]), .D (nx40390), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40391 (.Y (nx40390), .A0 (ram_75__2), .A1 (nx65854), .S0 (nx64020
             )) ;
    dffr reg_ram_74__2 (.Q (ram_74__2), .QB (\$dummy [603]), .D (nx40400), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40401 (.Y (nx40400), .A0 (ram_74__2), .A1 (nx65856), .S0 (nx64024
             )) ;
    aoi22 ix57105 (.Y (nx57104), .A0 (ram_76__2), .A1 (nx64954), .B0 (ram_77__2)
          , .B1 (nx64992)) ;
    dffr reg_ram_76__2 (.Q (ram_76__2), .QB (\$dummy [604]), .D (nx40380), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40381 (.Y (nx40380), .A0 (ram_76__2), .A1 (nx65856), .S0 (nx64016
             )) ;
    dffr reg_ram_77__2 (.Q (ram_77__2), .QB (\$dummy [605]), .D (nx40370), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40371 (.Y (nx40370), .A0 (ram_77__2), .A1 (nx65856), .S0 (nx64012
             )) ;
    aoi22 ix57113 (.Y (nx57112), .A0 (ram_79__2), .A1 (nx65030), .B0 (ram_78__2)
          , .B1 (nx65068)) ;
    dffr reg_ram_79__2 (.Q (ram_79__2), .QB (\$dummy [606]), .D (nx40350), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40351 (.Y (nx40350), .A0 (ram_79__2), .A1 (nx65856), .S0 (nx64004
             )) ;
    dffr reg_ram_78__2 (.Q (ram_78__2), .QB (\$dummy [607]), .D (nx40360), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40361 (.Y (nx40360), .A0 (ram_78__2), .A1 (nx65856), .S0 (nx64008
             )) ;
    oai21 ix57121 (.Y (nx57120), .A0 (nx9046), .A1 (nx8968), .B0 (nx65120)) ;
    nand04 ix9047 (.Y (nx9046), .A0 (nx57123), .A1 (nx57131), .A2 (nx57139), .A3 (
           nx57147)) ;
    aoi22 ix57124 (.Y (nx57123), .A0 (ram_48__2), .A1 (nx64498), .B0 (ram_49__2)
          , .B1 (nx64536)) ;
    dffr reg_ram_48__2 (.Q (ram_48__2), .QB (\$dummy [608]), .D (nx40340), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40341 (.Y (nx40340), .A0 (ram_48__2), .A1 (nx65856), .S0 (nx63994
             )) ;
    dffr reg_ram_49__2 (.Q (ram_49__2), .QB (\$dummy [609]), .D (nx40330), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40331 (.Y (nx40330), .A0 (ram_49__2), .A1 (nx65856), .S0 (nx63990
             )) ;
    aoi22 ix57132 (.Y (nx57131), .A0 (ram_51__2), .A1 (nx64574), .B0 (ram_50__2)
          , .B1 (nx64612)) ;
    dffr reg_ram_51__2 (.Q (ram_51__2), .QB (\$dummy [610]), .D (nx40310), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40311 (.Y (nx40310), .A0 (ram_51__2), .A1 (nx65858), .S0 (nx63982
             )) ;
    dffr reg_ram_50__2 (.Q (ram_50__2), .QB (\$dummy [611]), .D (nx40320), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40321 (.Y (nx40320), .A0 (ram_50__2), .A1 (nx65858), .S0 (nx63986
             )) ;
    aoi22 ix57140 (.Y (nx57139), .A0 (ram_52__2), .A1 (nx64650), .B0 (ram_53__2)
          , .B1 (nx64688)) ;
    dffr reg_ram_52__2 (.Q (ram_52__2), .QB (\$dummy [612]), .D (nx40300), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40301 (.Y (nx40300), .A0 (ram_52__2), .A1 (nx65858), .S0 (nx63978
             )) ;
    dffr reg_ram_53__2 (.Q (ram_53__2), .QB (\$dummy [613]), .D (nx40290), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40291 (.Y (nx40290), .A0 (ram_53__2), .A1 (nx65858), .S0 (nx63974
             )) ;
    aoi22 ix57148 (.Y (nx57147), .A0 (ram_55__2), .A1 (nx64726), .B0 (ram_54__2)
          , .B1 (nx64764)) ;
    dffr reg_ram_55__2 (.Q (ram_55__2), .QB (\$dummy [614]), .D (nx40270), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40271 (.Y (nx40270), .A0 (ram_55__2), .A1 (nx65858), .S0 (nx63966
             )) ;
    dffr reg_ram_54__2 (.Q (ram_54__2), .QB (\$dummy [615]), .D (nx40280), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40281 (.Y (nx40280), .A0 (ram_54__2), .A1 (nx65858), .S0 (nx63970
             )) ;
    nand04 ix8969 (.Y (nx8968), .A0 (nx57156), .A1 (nx57164), .A2 (nx57172), .A3 (
           nx57180)) ;
    aoi22 ix57157 (.Y (nx57156), .A0 (ram_56__2), .A1 (nx64802), .B0 (ram_57__2)
          , .B1 (nx64840)) ;
    dffr reg_ram_56__2 (.Q (ram_56__2), .QB (\$dummy [616]), .D (nx40260), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40261 (.Y (nx40260), .A0 (ram_56__2), .A1 (nx65858), .S0 (nx63962
             )) ;
    dffr reg_ram_57__2 (.Q (ram_57__2), .QB (\$dummy [617]), .D (nx40250), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40251 (.Y (nx40250), .A0 (ram_57__2), .A1 (nx65860), .S0 (nx63958
             )) ;
    aoi22 ix57165 (.Y (nx57164), .A0 (ram_59__2), .A1 (nx64878), .B0 (ram_58__2)
          , .B1 (nx64916)) ;
    dffr reg_ram_59__2 (.Q (ram_59__2), .QB (\$dummy [618]), .D (nx40230), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40231 (.Y (nx40230), .A0 (ram_59__2), .A1 (nx65860), .S0 (nx63950
             )) ;
    dffr reg_ram_58__2 (.Q (ram_58__2), .QB (\$dummy [619]), .D (nx40240), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40241 (.Y (nx40240), .A0 (ram_58__2), .A1 (nx65860), .S0 (nx63954
             )) ;
    aoi22 ix57173 (.Y (nx57172), .A0 (ram_60__2), .A1 (nx64954), .B0 (ram_61__2)
          , .B1 (nx64992)) ;
    dffr reg_ram_60__2 (.Q (ram_60__2), .QB (\$dummy [620]), .D (nx40220), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40221 (.Y (nx40220), .A0 (ram_60__2), .A1 (nx65860), .S0 (nx63946
             )) ;
    dffr reg_ram_61__2 (.Q (ram_61__2), .QB (\$dummy [621]), .D (nx40210), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40211 (.Y (nx40210), .A0 (ram_61__2), .A1 (nx65860), .S0 (nx63942
             )) ;
    aoi22 ix57181 (.Y (nx57180), .A0 (ram_63__2), .A1 (nx65030), .B0 (ram_62__2)
          , .B1 (nx65068)) ;
    dffr reg_ram_63__2 (.Q (ram_63__2), .QB (\$dummy [622]), .D (nx40190), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40191 (.Y (nx40190), .A0 (ram_63__2), .A1 (nx65860), .S0 (nx63934
             )) ;
    dffr reg_ram_62__2 (.Q (ram_62__2), .QB (\$dummy [623]), .D (nx40200), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40201 (.Y (nx40200), .A0 (ram_62__2), .A1 (nx65860), .S0 (nx63938
             )) ;
    oai21 ix57189 (.Y (nx57188), .A0 (nx8884), .A1 (nx8806), .B0 (nx65124)) ;
    nand04 ix8885 (.Y (nx8884), .A0 (nx57191), .A1 (nx57199), .A2 (nx57207), .A3 (
           nx57215)) ;
    aoi22 ix57192 (.Y (nx57191), .A0 (ram_32__2), .A1 (nx64498), .B0 (ram_33__2)
          , .B1 (nx64536)) ;
    dffr reg_ram_32__2 (.Q (ram_32__2), .QB (\$dummy [624]), .D (nx40180), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40181 (.Y (nx40180), .A0 (ram_32__2), .A1 (nx65862), .S0 (nx63924
             )) ;
    dffr reg_ram_33__2 (.Q (ram_33__2), .QB (\$dummy [625]), .D (nx40170), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40171 (.Y (nx40170), .A0 (ram_33__2), .A1 (nx65862), .S0 (nx63920
             )) ;
    aoi22 ix57200 (.Y (nx57199), .A0 (ram_35__2), .A1 (nx64574), .B0 (ram_34__2)
          , .B1 (nx64612)) ;
    dffr reg_ram_35__2 (.Q (ram_35__2), .QB (\$dummy [626]), .D (nx40150), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40151 (.Y (nx40150), .A0 (ram_35__2), .A1 (nx65862), .S0 (nx63912
             )) ;
    dffr reg_ram_34__2 (.Q (ram_34__2), .QB (\$dummy [627]), .D (nx40160), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40161 (.Y (nx40160), .A0 (ram_34__2), .A1 (nx65862), .S0 (nx63916
             )) ;
    aoi22 ix57208 (.Y (nx57207), .A0 (ram_36__2), .A1 (nx64650), .B0 (ram_37__2)
          , .B1 (nx64688)) ;
    dffr reg_ram_36__2 (.Q (ram_36__2), .QB (\$dummy [628]), .D (nx40140), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40141 (.Y (nx40140), .A0 (ram_36__2), .A1 (nx65862), .S0 (nx63908
             )) ;
    dffr reg_ram_37__2 (.Q (ram_37__2), .QB (\$dummy [629]), .D (nx40130), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40131 (.Y (nx40130), .A0 (ram_37__2), .A1 (nx65862), .S0 (nx63904
             )) ;
    aoi22 ix57216 (.Y (nx57215), .A0 (ram_39__2), .A1 (nx64726), .B0 (ram_38__2)
          , .B1 (nx64764)) ;
    dffr reg_ram_39__2 (.Q (ram_39__2), .QB (\$dummy [630]), .D (nx40110), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40111 (.Y (nx40110), .A0 (ram_39__2), .A1 (nx65862), .S0 (nx63896
             )) ;
    dffr reg_ram_38__2 (.Q (ram_38__2), .QB (\$dummy [631]), .D (nx40120), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40121 (.Y (nx40120), .A0 (ram_38__2), .A1 (nx65864), .S0 (nx63900
             )) ;
    nand04 ix8807 (.Y (nx8806), .A0 (nx57224), .A1 (nx57232), .A2 (nx57240), .A3 (
           nx57248)) ;
    aoi22 ix57225 (.Y (nx57224), .A0 (ram_40__2), .A1 (nx64802), .B0 (ram_41__2)
          , .B1 (nx64840)) ;
    dffr reg_ram_40__2 (.Q (ram_40__2), .QB (\$dummy [632]), .D (nx40100), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40101 (.Y (nx40100), .A0 (ram_40__2), .A1 (nx65864), .S0 (nx63892
             )) ;
    dffr reg_ram_41__2 (.Q (ram_41__2), .QB (\$dummy [633]), .D (nx40090), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40091 (.Y (nx40090), .A0 (ram_41__2), .A1 (nx65864), .S0 (nx63888
             )) ;
    aoi22 ix57233 (.Y (nx57232), .A0 (ram_43__2), .A1 (nx64878), .B0 (ram_42__2)
          , .B1 (nx64916)) ;
    dffr reg_ram_43__2 (.Q (ram_43__2), .QB (\$dummy [634]), .D (nx40070), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40071 (.Y (nx40070), .A0 (ram_43__2), .A1 (nx65864), .S0 (nx63880
             )) ;
    dffr reg_ram_42__2 (.Q (ram_42__2), .QB (\$dummy [635]), .D (nx40080), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40081 (.Y (nx40080), .A0 (ram_42__2), .A1 (nx65864), .S0 (nx63884
             )) ;
    aoi22 ix57241 (.Y (nx57240), .A0 (ram_44__2), .A1 (nx64954), .B0 (ram_45__2)
          , .B1 (nx64992)) ;
    dffr reg_ram_44__2 (.Q (ram_44__2), .QB (\$dummy [636]), .D (nx40060), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40061 (.Y (nx40060), .A0 (ram_44__2), .A1 (nx65864), .S0 (nx63876
             )) ;
    dffr reg_ram_45__2 (.Q (ram_45__2), .QB (\$dummy [637]), .D (nx40050), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40051 (.Y (nx40050), .A0 (ram_45__2), .A1 (nx65864), .S0 (nx63872
             )) ;
    aoi22 ix57249 (.Y (nx57248), .A0 (ram_47__2), .A1 (nx65030), .B0 (ram_46__2)
          , .B1 (nx65068)) ;
    dffr reg_ram_47__2 (.Q (ram_47__2), .QB (\$dummy [638]), .D (nx40030), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40031 (.Y (nx40030), .A0 (ram_47__2), .A1 (nx65866), .S0 (nx63864
             )) ;
    dffr reg_ram_46__2 (.Q (ram_46__2), .QB (\$dummy [639]), .D (nx40040), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40041 (.Y (nx40040), .A0 (ram_46__2), .A1 (nx65866), .S0 (nx63868
             )) ;
    nand04 ix8727 (.Y (nx8726), .A0 (nx57257), .A1 (nx57325), .A2 (nx57393), .A3 (
           nx57461)) ;
    oai21 ix57258 (.Y (nx57257), .A0 (nx8716), .A1 (nx8638), .B0 (nx65128)) ;
    nand04 ix8717 (.Y (nx8716), .A0 (nx57260), .A1 (nx57268), .A2 (nx57276), .A3 (
           nx57284)) ;
    aoi22 ix57261 (.Y (nx57260), .A0 (ram_16__2), .A1 (nx64498), .B0 (ram_17__2)
          , .B1 (nx64536)) ;
    dffr reg_ram_16__2 (.Q (ram_16__2), .QB (\$dummy [640]), .D (nx40020), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40021 (.Y (nx40020), .A0 (ram_16__2), .A1 (nx65866), .S0 (nx63854
             )) ;
    dffr reg_ram_17__2 (.Q (ram_17__2), .QB (\$dummy [641]), .D (nx40010), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40011 (.Y (nx40010), .A0 (ram_17__2), .A1 (nx65866), .S0 (nx63850
             )) ;
    aoi22 ix57269 (.Y (nx57268), .A0 (ram_19__2), .A1 (nx64574), .B0 (ram_18__2)
          , .B1 (nx64612)) ;
    dffr reg_ram_19__2 (.Q (ram_19__2), .QB (\$dummy [642]), .D (nx39990), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39991 (.Y (nx39990), .A0 (ram_19__2), .A1 (nx65866), .S0 (nx63842
             )) ;
    dffr reg_ram_18__2 (.Q (ram_18__2), .QB (\$dummy [643]), .D (nx40000), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix40001 (.Y (nx40000), .A0 (ram_18__2), .A1 (nx65866), .S0 (nx63846
             )) ;
    aoi22 ix57277 (.Y (nx57276), .A0 (ram_20__2), .A1 (nx64650), .B0 (ram_21__2)
          , .B1 (nx64688)) ;
    dffr reg_ram_20__2 (.Q (ram_20__2), .QB (\$dummy [644]), .D (nx39980), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39981 (.Y (nx39980), .A0 (ram_20__2), .A1 (nx65866), .S0 (nx63838
             )) ;
    dffr reg_ram_21__2 (.Q (ram_21__2), .QB (\$dummy [645]), .D (nx39970), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39971 (.Y (nx39970), .A0 (ram_21__2), .A1 (nx65868), .S0 (nx63834
             )) ;
    aoi22 ix57285 (.Y (nx57284), .A0 (ram_23__2), .A1 (nx64726), .B0 (ram_22__2)
          , .B1 (nx64764)) ;
    dffr reg_ram_23__2 (.Q (ram_23__2), .QB (\$dummy [646]), .D (nx39950), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39951 (.Y (nx39950), .A0 (ram_23__2), .A1 (nx65868), .S0 (nx63826
             )) ;
    dffr reg_ram_22__2 (.Q (ram_22__2), .QB (\$dummy [647]), .D (nx39960), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39961 (.Y (nx39960), .A0 (ram_22__2), .A1 (nx65868), .S0 (nx63830
             )) ;
    nand04 ix8639 (.Y (nx8638), .A0 (nx57293), .A1 (nx57301), .A2 (nx57309), .A3 (
           nx57317)) ;
    aoi22 ix57294 (.Y (nx57293), .A0 (ram_24__2), .A1 (nx64802), .B0 (ram_25__2)
          , .B1 (nx64840)) ;
    dffr reg_ram_24__2 (.Q (ram_24__2), .QB (\$dummy [648]), .D (nx39940), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39941 (.Y (nx39940), .A0 (ram_24__2), .A1 (nx65868), .S0 (nx63822
             )) ;
    dffr reg_ram_25__2 (.Q (ram_25__2), .QB (\$dummy [649]), .D (nx39930), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39931 (.Y (nx39930), .A0 (ram_25__2), .A1 (nx65868), .S0 (nx63818
             )) ;
    aoi22 ix57302 (.Y (nx57301), .A0 (ram_27__2), .A1 (nx64878), .B0 (ram_26__2)
          , .B1 (nx64916)) ;
    dffr reg_ram_27__2 (.Q (ram_27__2), .QB (\$dummy [650]), .D (nx39910), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39911 (.Y (nx39910), .A0 (ram_27__2), .A1 (nx65868), .S0 (nx63810
             )) ;
    dffr reg_ram_26__2 (.Q (ram_26__2), .QB (\$dummy [651]), .D (nx39920), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39921 (.Y (nx39920), .A0 (ram_26__2), .A1 (nx65868), .S0 (nx63814
             )) ;
    aoi22 ix57310 (.Y (nx57309), .A0 (ram_28__2), .A1 (nx64954), .B0 (ram_29__2)
          , .B1 (nx64992)) ;
    dffr reg_ram_28__2 (.Q (ram_28__2), .QB (\$dummy [652]), .D (nx39900), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39901 (.Y (nx39900), .A0 (ram_28__2), .A1 (nx65870), .S0 (nx63806
             )) ;
    dffr reg_ram_29__2 (.Q (ram_29__2), .QB (\$dummy [653]), .D (nx39890), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39891 (.Y (nx39890), .A0 (ram_29__2), .A1 (nx65870), .S0 (nx63802
             )) ;
    aoi22 ix57318 (.Y (nx57317), .A0 (ram_31__2), .A1 (nx65030), .B0 (ram_30__2)
          , .B1 (nx65068)) ;
    dffr reg_ram_31__2 (.Q (ram_31__2), .QB (\$dummy [654]), .D (nx39870), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39871 (.Y (nx39870), .A0 (ram_31__2), .A1 (nx65870), .S0 (nx63794
             )) ;
    dffr reg_ram_30__2 (.Q (ram_30__2), .QB (\$dummy [655]), .D (nx39880), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39881 (.Y (nx39880), .A0 (ram_30__2), .A1 (nx65870), .S0 (nx63798
             )) ;
    oai21 ix57326 (.Y (nx57325), .A0 (nx8554), .A1 (nx8476), .B0 (nx65142)) ;
    nand04 ix8555 (.Y (nx8554), .A0 (nx57328), .A1 (nx57336), .A2 (nx57344), .A3 (
           nx57352)) ;
    aoi22 ix57329 (.Y (nx57328), .A0 (ram_0__2), .A1 (nx64500), .B0 (ram_1__2), 
          .B1 (nx64538)) ;
    dffr reg_ram_0__2 (.Q (ram_0__2), .QB (\$dummy [656]), .D (nx39860), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39861 (.Y (nx39860), .A0 (nx65870), .A1 (ram_0__2), .S0 (nx65132)
             ) ;
    dffr reg_ram_1__2 (.Q (ram_1__2), .QB (\$dummy [657]), .D (nx39850), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39851 (.Y (nx39850), .A0 (nx65870), .A1 (ram_1__2), .S0 (nx65146)
             ) ;
    aoi22 ix57337 (.Y (nx57336), .A0 (ram_3__2), .A1 (nx64576), .B0 (ram_2__2), 
          .B1 (nx64614)) ;
    dffr reg_ram_3__2 (.Q (ram_3__2), .QB (\$dummy [658]), .D (nx39830), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39831 (.Y (nx39830), .A0 (nx65870), .A1 (ram_3__2), .S0 (nx65150)
             ) ;
    dffr reg_ram_2__2 (.Q (ram_2__2), .QB (\$dummy [659]), .D (nx39840), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39841 (.Y (nx39840), .A0 (nx65872), .A1 (ram_2__2), .S0 (nx65154)
             ) ;
    aoi22 ix57345 (.Y (nx57344), .A0 (ram_4__2), .A1 (nx64652), .B0 (ram_5__2), 
          .B1 (nx64690)) ;
    dffr reg_ram_4__2 (.Q (ram_4__2), .QB (\$dummy [660]), .D (nx39820), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39821 (.Y (nx39820), .A0 (nx65872), .A1 (ram_4__2), .S0 (nx65158)
             ) ;
    dffr reg_ram_5__2 (.Q (ram_5__2), .QB (\$dummy [661]), .D (nx39810), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39811 (.Y (nx39810), .A0 (nx65872), .A1 (ram_5__2), .S0 (nx65162)
             ) ;
    aoi22 ix57353 (.Y (nx57352), .A0 (ram_7__2), .A1 (nx64728), .B0 (ram_6__2), 
          .B1 (nx64766)) ;
    dffr reg_ram_7__2 (.Q (ram_7__2), .QB (\$dummy [662]), .D (nx39790), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39791 (.Y (nx39790), .A0 (nx65872), .A1 (ram_7__2), .S0 (nx65166)
             ) ;
    dffr reg_ram_6__2 (.Q (ram_6__2), .QB (\$dummy [663]), .D (nx39800), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39801 (.Y (nx39800), .A0 (nx65872), .A1 (ram_6__2), .S0 (nx65170)
             ) ;
    nand04 ix8477 (.Y (nx8476), .A0 (nx57361), .A1 (nx57369), .A2 (nx57377), .A3 (
           nx57385)) ;
    aoi22 ix57362 (.Y (nx57361), .A0 (ram_8__2), .A1 (nx64804), .B0 (ram_9__2), 
          .B1 (nx64842)) ;
    dffr reg_ram_8__2 (.Q (ram_8__2), .QB (\$dummy [664]), .D (nx39780), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39781 (.Y (nx39780), .A0 (nx65872), .A1 (ram_8__2), .S0 (nx65174)
             ) ;
    dffr reg_ram_9__2 (.Q (ram_9__2), .QB (\$dummy [665]), .D (nx39770), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39771 (.Y (nx39770), .A0 (nx65872), .A1 (ram_9__2), .S0 (nx65178)
             ) ;
    aoi22 ix57370 (.Y (nx57369), .A0 (ram_11__2), .A1 (nx64880), .B0 (ram_10__2)
          , .B1 (nx64918)) ;
    dffr reg_ram_11__2 (.Q (ram_11__2), .QB (\$dummy [666]), .D (nx39750), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39751 (.Y (nx39750), .A0 (nx65874), .A1 (ram_11__2), .S0 (nx65182
             )) ;
    dffr reg_ram_10__2 (.Q (ram_10__2), .QB (\$dummy [667]), .D (nx39760), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39761 (.Y (nx39760), .A0 (nx65874), .A1 (ram_10__2), .S0 (nx65186
             )) ;
    aoi22 ix57378 (.Y (nx57377), .A0 (ram_12__2), .A1 (nx64956), .B0 (ram_13__2)
          , .B1 (nx64994)) ;
    dffr reg_ram_12__2 (.Q (ram_12__2), .QB (\$dummy [668]), .D (nx39740), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39741 (.Y (nx39740), .A0 (nx65874), .A1 (ram_12__2), .S0 (nx65190
             )) ;
    dffr reg_ram_13__2 (.Q (ram_13__2), .QB (\$dummy [669]), .D (nx39730), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39731 (.Y (nx39730), .A0 (nx65874), .A1 (ram_13__2), .S0 (nx65194
             )) ;
    aoi22 ix57386 (.Y (nx57385), .A0 (ram_15__2), .A1 (nx65032), .B0 (ram_14__2)
          , .B1 (nx65070)) ;
    dffr reg_ram_15__2 (.Q (ram_15__2), .QB (\$dummy [670]), .D (nx39710), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39711 (.Y (nx39710), .A0 (nx65874), .A1 (ram_15__2), .S0 (nx65198
             )) ;
    dffr reg_ram_14__2 (.Q (ram_14__2), .QB (\$dummy [671]), .D (nx39720), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39721 (.Y (nx39720), .A0 (nx65874), .A1 (ram_14__2), .S0 (nx65202
             )) ;
    oai21 ix57394 (.Y (nx57393), .A0 (nx8390), .A1 (nx8312), .B0 (nx65206)) ;
    nand04 ix8391 (.Y (nx8390), .A0 (nx57396), .A1 (nx57404), .A2 (nx57412), .A3 (
           nx57420)) ;
    aoi22 ix57397 (.Y (nx57396), .A0 (ram_96__2), .A1 (nx64500), .B0 (ram_97__2)
          , .B1 (nx64538)) ;
    dffr reg_ram_96__2 (.Q (ram_96__2), .QB (\$dummy [672]), .D (nx39700), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39701 (.Y (nx39700), .A0 (ram_96__2), .A1 (nx65874), .S0 (nx63784
             )) ;
    dffr reg_ram_97__2 (.Q (ram_97__2), .QB (\$dummy [673]), .D (nx39690), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39691 (.Y (nx39690), .A0 (ram_97__2), .A1 (nx65876), .S0 (nx63780
             )) ;
    aoi22 ix57405 (.Y (nx57404), .A0 (ram_99__2), .A1 (nx64576), .B0 (ram_98__2)
          , .B1 (nx64614)) ;
    dffr reg_ram_99__2 (.Q (ram_99__2), .QB (\$dummy [674]), .D (nx39670), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39671 (.Y (nx39670), .A0 (ram_99__2), .A1 (nx65876), .S0 (nx63772
             )) ;
    dffr reg_ram_98__2 (.Q (ram_98__2), .QB (\$dummy [675]), .D (nx39680), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39681 (.Y (nx39680), .A0 (ram_98__2), .A1 (nx65876), .S0 (nx63776
             )) ;
    aoi22 ix57413 (.Y (nx57412), .A0 (ram_100__2), .A1 (nx64652), .B0 (
          ram_101__2), .B1 (nx64690)) ;
    dffr reg_ram_100__2 (.Q (ram_100__2), .QB (\$dummy [676]), .D (nx39660), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39661 (.Y (nx39660), .A0 (ram_100__2), .A1 (nx65876), .S0 (
             nx63768)) ;
    dffr reg_ram_101__2 (.Q (ram_101__2), .QB (\$dummy [677]), .D (nx39650), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39651 (.Y (nx39650), .A0 (ram_101__2), .A1 (nx65876), .S0 (
             nx63764)) ;
    aoi22 ix57421 (.Y (nx57420), .A0 (ram_103__2), .A1 (nx64728), .B0 (
          ram_102__2), .B1 (nx64766)) ;
    dffr reg_ram_103__2 (.Q (ram_103__2), .QB (\$dummy [678]), .D (nx39630), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39631 (.Y (nx39630), .A0 (ram_103__2), .A1 (nx65876), .S0 (
             nx63756)) ;
    dffr reg_ram_102__2 (.Q (ram_102__2), .QB (\$dummy [679]), .D (nx39640), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39641 (.Y (nx39640), .A0 (ram_102__2), .A1 (nx65876), .S0 (
             nx63760)) ;
    nand04 ix8313 (.Y (nx8312), .A0 (nx57429), .A1 (nx57437), .A2 (nx57445), .A3 (
           nx57453)) ;
    aoi22 ix57430 (.Y (nx57429), .A0 (ram_104__2), .A1 (nx64804), .B0 (
          ram_105__2), .B1 (nx64842)) ;
    dffr reg_ram_104__2 (.Q (ram_104__2), .QB (\$dummy [680]), .D (nx39620), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39621 (.Y (nx39620), .A0 (ram_104__2), .A1 (nx65878), .S0 (
             nx63752)) ;
    dffr reg_ram_105__2 (.Q (ram_105__2), .QB (\$dummy [681]), .D (nx39610), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39611 (.Y (nx39610), .A0 (ram_105__2), .A1 (nx65878), .S0 (
             nx63748)) ;
    aoi22 ix57438 (.Y (nx57437), .A0 (ram_107__2), .A1 (nx64880), .B0 (
          ram_106__2), .B1 (nx64918)) ;
    dffr reg_ram_107__2 (.Q (ram_107__2), .QB (\$dummy [682]), .D (nx39590), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39591 (.Y (nx39590), .A0 (ram_107__2), .A1 (nx65878), .S0 (
             nx63740)) ;
    dffr reg_ram_106__2 (.Q (ram_106__2), .QB (\$dummy [683]), .D (nx39600), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39601 (.Y (nx39600), .A0 (ram_106__2), .A1 (nx65878), .S0 (
             nx63744)) ;
    aoi22 ix57446 (.Y (nx57445), .A0 (ram_108__2), .A1 (nx64956), .B0 (
          ram_109__2), .B1 (nx64994)) ;
    dffr reg_ram_108__2 (.Q (ram_108__2), .QB (\$dummy [684]), .D (nx39580), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39581 (.Y (nx39580), .A0 (ram_108__2), .A1 (nx65878), .S0 (
             nx63736)) ;
    dffr reg_ram_109__2 (.Q (ram_109__2), .QB (\$dummy [685]), .D (nx39570), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39571 (.Y (nx39570), .A0 (ram_109__2), .A1 (nx65878), .S0 (
             nx63732)) ;
    aoi22 ix57454 (.Y (nx57453), .A0 (ram_111__2), .A1 (nx65032), .B0 (
          ram_110__2), .B1 (nx65070)) ;
    dffr reg_ram_111__2 (.Q (ram_111__2), .QB (\$dummy [686]), .D (nx39550), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39551 (.Y (nx39550), .A0 (ram_111__2), .A1 (nx65878), .S0 (
             nx63724)) ;
    dffr reg_ram_110__2 (.Q (ram_110__2), .QB (\$dummy [687]), .D (nx39560), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39561 (.Y (nx39560), .A0 (ram_110__2), .A1 (nx65880), .S0 (
             nx63728)) ;
    oai21 ix57462 (.Y (nx57461), .A0 (nx8228), .A1 (nx8150), .B0 (nx65210)) ;
    nand04 ix8229 (.Y (nx8228), .A0 (nx57464), .A1 (nx57472), .A2 (nx57480), .A3 (
           nx57488)) ;
    aoi22 ix57465 (.Y (nx57464), .A0 (ram_112__2), .A1 (nx64500), .B0 (
          ram_113__2), .B1 (nx64538)) ;
    dffr reg_ram_112__2 (.Q (ram_112__2), .QB (\$dummy [688]), .D (nx39540), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39541 (.Y (nx39540), .A0 (ram_112__2), .A1 (nx65880), .S0 (
             nx63714)) ;
    dffr reg_ram_113__2 (.Q (ram_113__2), .QB (\$dummy [689]), .D (nx39530), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39531 (.Y (nx39530), .A0 (ram_113__2), .A1 (nx65880), .S0 (
             nx63710)) ;
    aoi22 ix57473 (.Y (nx57472), .A0 (ram_115__2), .A1 (nx64576), .B0 (
          ram_114__2), .B1 (nx64614)) ;
    dffr reg_ram_115__2 (.Q (ram_115__2), .QB (\$dummy [690]), .D (nx39510), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39511 (.Y (nx39510), .A0 (ram_115__2), .A1 (nx65880), .S0 (
             nx63702)) ;
    dffr reg_ram_114__2 (.Q (ram_114__2), .QB (\$dummy [691]), .D (nx39520), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39521 (.Y (nx39520), .A0 (ram_114__2), .A1 (nx65880), .S0 (
             nx63706)) ;
    aoi22 ix57481 (.Y (nx57480), .A0 (ram_116__2), .A1 (nx64652), .B0 (
          ram_117__2), .B1 (nx64690)) ;
    dffr reg_ram_116__2 (.Q (ram_116__2), .QB (\$dummy [692]), .D (nx39500), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39501 (.Y (nx39500), .A0 (ram_116__2), .A1 (nx65880), .S0 (
             nx63698)) ;
    dffr reg_ram_117__2 (.Q (ram_117__2), .QB (\$dummy [693]), .D (nx39490), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39491 (.Y (nx39490), .A0 (ram_117__2), .A1 (nx65880), .S0 (
             nx63694)) ;
    aoi22 ix57489 (.Y (nx57488), .A0 (ram_119__2), .A1 (nx64728), .B0 (
          ram_118__2), .B1 (nx64766)) ;
    dffr reg_ram_119__2 (.Q (ram_119__2), .QB (\$dummy [694]), .D (nx39470), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39471 (.Y (nx39470), .A0 (ram_119__2), .A1 (nx65882), .S0 (
             nx63686)) ;
    dffr reg_ram_118__2 (.Q (ram_118__2), .QB (\$dummy [695]), .D (nx39480), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39481 (.Y (nx39480), .A0 (ram_118__2), .A1 (nx65882), .S0 (
             nx63690)) ;
    nand04 ix8151 (.Y (nx8150), .A0 (nx57497), .A1 (nx57505), .A2 (nx57513), .A3 (
           nx57521)) ;
    aoi22 ix57498 (.Y (nx57497), .A0 (ram_120__2), .A1 (nx64804), .B0 (
          ram_121__2), .B1 (nx64842)) ;
    dffr reg_ram_120__2 (.Q (ram_120__2), .QB (\$dummy [696]), .D (nx39460), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39461 (.Y (nx39460), .A0 (ram_120__2), .A1 (nx65882), .S0 (
             nx63682)) ;
    dffr reg_ram_121__2 (.Q (ram_121__2), .QB (\$dummy [697]), .D (nx39450), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39451 (.Y (nx39450), .A0 (ram_121__2), .A1 (nx65882), .S0 (
             nx63678)) ;
    aoi22 ix57506 (.Y (nx57505), .A0 (ram_123__2), .A1 (nx64880), .B0 (
          ram_122__2), .B1 (nx64918)) ;
    dffr reg_ram_123__2 (.Q (ram_123__2), .QB (\$dummy [698]), .D (nx39430), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39431 (.Y (nx39430), .A0 (ram_123__2), .A1 (nx65882), .S0 (
             nx63670)) ;
    dffr reg_ram_122__2 (.Q (ram_122__2), .QB (\$dummy [699]), .D (nx39440), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39441 (.Y (nx39440), .A0 (ram_122__2), .A1 (nx65882), .S0 (
             nx63674)) ;
    aoi22 ix57514 (.Y (nx57513), .A0 (ram_124__2), .A1 (nx64956), .B0 (
          ram_125__2), .B1 (nx64994)) ;
    dffr reg_ram_124__2 (.Q (ram_124__2), .QB (\$dummy [700]), .D (nx39420), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39421 (.Y (nx39420), .A0 (ram_124__2), .A1 (nx65882), .S0 (
             nx63666)) ;
    dffr reg_ram_125__2 (.Q (ram_125__2), .QB (\$dummy [701]), .D (nx39410), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39411 (.Y (nx39410), .A0 (ram_125__2), .A1 (nx65884), .S0 (
             nx63662)) ;
    aoi22 ix57522 (.Y (nx57521), .A0 (ram_127__2), .A1 (nx65032), .B0 (
          ram_126__2), .B1 (nx65070)) ;
    dffr reg_ram_127__2 (.Q (ram_127__2), .QB (\$dummy [702]), .D (nx39390), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39391 (.Y (nx39390), .A0 (ram_127__2), .A1 (nx65884), .S0 (
             nx63654)) ;
    dffr reg_ram_126__2 (.Q (ram_126__2), .QB (\$dummy [703]), .D (nx39400), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39401 (.Y (nx39400), .A0 (ram_126__2), .A1 (nx65884), .S0 (
             nx63658)) ;
    nand04 ix8073 (.Y (nx8072), .A0 (nx57530), .A1 (nx57598), .A2 (nx57666), .A3 (
           nx57734)) ;
    oai21 ix57531 (.Y (nx57530), .A0 (nx8062), .A1 (nx7984), .B0 (nx65214)) ;
    nand04 ix8063 (.Y (nx8062), .A0 (nx57533), .A1 (nx57541), .A2 (nx57549), .A3 (
           nx57557)) ;
    aoi22 ix57534 (.Y (nx57533), .A0 (ram_128__2), .A1 (nx64500), .B0 (
          ram_129__2), .B1 (nx64538)) ;
    dffr reg_ram_128__2 (.Q (ram_128__2), .QB (\$dummy [704]), .D (nx39380), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39381 (.Y (nx39380), .A0 (ram_128__2), .A1 (nx65884), .S0 (
             nx63644)) ;
    dffr reg_ram_129__2 (.Q (ram_129__2), .QB (\$dummy [705]), .D (nx39370), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39371 (.Y (nx39370), .A0 (ram_129__2), .A1 (nx65884), .S0 (
             nx63640)) ;
    aoi22 ix57542 (.Y (nx57541), .A0 (ram_131__2), .A1 (nx64576), .B0 (
          ram_130__2), .B1 (nx64614)) ;
    dffr reg_ram_131__2 (.Q (ram_131__2), .QB (\$dummy [706]), .D (nx39350), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39351 (.Y (nx39350), .A0 (ram_131__2), .A1 (nx65884), .S0 (
             nx63632)) ;
    dffr reg_ram_130__2 (.Q (ram_130__2), .QB (\$dummy [707]), .D (nx39360), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39361 (.Y (nx39360), .A0 (ram_130__2), .A1 (nx65884), .S0 (
             nx63636)) ;
    aoi22 ix57550 (.Y (nx57549), .A0 (ram_132__2), .A1 (nx64652), .B0 (
          ram_133__2), .B1 (nx64690)) ;
    dffr reg_ram_132__2 (.Q (ram_132__2), .QB (\$dummy [708]), .D (nx39340), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39341 (.Y (nx39340), .A0 (ram_132__2), .A1 (nx65886), .S0 (
             nx63628)) ;
    dffr reg_ram_133__2 (.Q (ram_133__2), .QB (\$dummy [709]), .D (nx39330), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39331 (.Y (nx39330), .A0 (ram_133__2), .A1 (nx65886), .S0 (
             nx63624)) ;
    aoi22 ix57558 (.Y (nx57557), .A0 (ram_135__2), .A1 (nx64728), .B0 (
          ram_134__2), .B1 (nx64766)) ;
    dffr reg_ram_135__2 (.Q (ram_135__2), .QB (\$dummy [710]), .D (nx39310), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39311 (.Y (nx39310), .A0 (ram_135__2), .A1 (nx65886), .S0 (
             nx63616)) ;
    dffr reg_ram_134__2 (.Q (ram_134__2), .QB (\$dummy [711]), .D (nx39320), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39321 (.Y (nx39320), .A0 (ram_134__2), .A1 (nx65886), .S0 (
             nx63620)) ;
    nand04 ix7985 (.Y (nx7984), .A0 (nx57566), .A1 (nx57574), .A2 (nx57582), .A3 (
           nx57590)) ;
    aoi22 ix57567 (.Y (nx57566), .A0 (ram_136__2), .A1 (nx64804), .B0 (
          ram_137__2), .B1 (nx64842)) ;
    dffr reg_ram_136__2 (.Q (ram_136__2), .QB (\$dummy [712]), .D (nx39300), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39301 (.Y (nx39300), .A0 (ram_136__2), .A1 (nx65886), .S0 (
             nx63612)) ;
    dffr reg_ram_137__2 (.Q (ram_137__2), .QB (\$dummy [713]), .D (nx39290), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39291 (.Y (nx39290), .A0 (ram_137__2), .A1 (nx65886), .S0 (
             nx63608)) ;
    aoi22 ix57575 (.Y (nx57574), .A0 (ram_139__2), .A1 (nx64880), .B0 (
          ram_138__2), .B1 (nx64918)) ;
    dffr reg_ram_139__2 (.Q (ram_139__2), .QB (\$dummy [714]), .D (nx39270), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39271 (.Y (nx39270), .A0 (ram_139__2), .A1 (nx65886), .S0 (
             nx63600)) ;
    dffr reg_ram_138__2 (.Q (ram_138__2), .QB (\$dummy [715]), .D (nx39280), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39281 (.Y (nx39280), .A0 (ram_138__2), .A1 (nx65888), .S0 (
             nx63604)) ;
    aoi22 ix57583 (.Y (nx57582), .A0 (ram_140__2), .A1 (nx64956), .B0 (
          ram_141__2), .B1 (nx64994)) ;
    dffr reg_ram_140__2 (.Q (ram_140__2), .QB (\$dummy [716]), .D (nx39260), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39261 (.Y (nx39260), .A0 (ram_140__2), .A1 (nx65888), .S0 (
             nx63596)) ;
    dffr reg_ram_141__2 (.Q (ram_141__2), .QB (\$dummy [717]), .D (nx39250), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39251 (.Y (nx39250), .A0 (ram_141__2), .A1 (nx65888), .S0 (
             nx63592)) ;
    aoi22 ix57591 (.Y (nx57590), .A0 (ram_143__2), .A1 (nx65032), .B0 (
          ram_142__2), .B1 (nx65070)) ;
    dffr reg_ram_143__2 (.Q (ram_143__2), .QB (\$dummy [718]), .D (nx39230), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39231 (.Y (nx39230), .A0 (ram_143__2), .A1 (nx65888), .S0 (
             nx63584)) ;
    dffr reg_ram_142__2 (.Q (ram_142__2), .QB (\$dummy [719]), .D (nx39240), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39241 (.Y (nx39240), .A0 (ram_142__2), .A1 (nx65888), .S0 (
             nx63588)) ;
    oai21 ix57599 (.Y (nx57598), .A0 (nx7900), .A1 (nx7822), .B0 (nx65218)) ;
    nand04 ix7901 (.Y (nx7900), .A0 (nx57601), .A1 (nx57609), .A2 (nx57617), .A3 (
           nx57625)) ;
    aoi22 ix57602 (.Y (nx57601), .A0 (ram_144__2), .A1 (nx64500), .B0 (
          ram_145__2), .B1 (nx64538)) ;
    dffr reg_ram_144__2 (.Q (ram_144__2), .QB (\$dummy [720]), .D (nx39220), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39221 (.Y (nx39220), .A0 (ram_144__2), .A1 (nx65888), .S0 (
             nx63574)) ;
    dffr reg_ram_145__2 (.Q (ram_145__2), .QB (\$dummy [721]), .D (nx39210), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39211 (.Y (nx39210), .A0 (ram_145__2), .A1 (nx65888), .S0 (
             nx63570)) ;
    aoi22 ix57610 (.Y (nx57609), .A0 (ram_147__2), .A1 (nx64576), .B0 (
          ram_146__2), .B1 (nx64614)) ;
    dffr reg_ram_147__2 (.Q (ram_147__2), .QB (\$dummy [722]), .D (nx39190), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39191 (.Y (nx39190), .A0 (ram_147__2), .A1 (nx65890), .S0 (
             nx63562)) ;
    dffr reg_ram_146__2 (.Q (ram_146__2), .QB (\$dummy [723]), .D (nx39200), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39201 (.Y (nx39200), .A0 (ram_146__2), .A1 (nx65890), .S0 (
             nx63566)) ;
    aoi22 ix57618 (.Y (nx57617), .A0 (ram_148__2), .A1 (nx64652), .B0 (
          ram_149__2), .B1 (nx64690)) ;
    dffr reg_ram_148__2 (.Q (ram_148__2), .QB (\$dummy [724]), .D (nx39180), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39181 (.Y (nx39180), .A0 (ram_148__2), .A1 (nx65890), .S0 (
             nx63558)) ;
    dffr reg_ram_149__2 (.Q (ram_149__2), .QB (\$dummy [725]), .D (nx39170), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39171 (.Y (nx39170), .A0 (ram_149__2), .A1 (nx65890), .S0 (
             nx63554)) ;
    aoi22 ix57626 (.Y (nx57625), .A0 (ram_151__2), .A1 (nx64728), .B0 (
          ram_150__2), .B1 (nx64766)) ;
    dffr reg_ram_151__2 (.Q (ram_151__2), .QB (\$dummy [726]), .D (nx39150), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39151 (.Y (nx39150), .A0 (ram_151__2), .A1 (nx65890), .S0 (
             nx63546)) ;
    dffr reg_ram_150__2 (.Q (ram_150__2), .QB (\$dummy [727]), .D (nx39160), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39161 (.Y (nx39160), .A0 (ram_150__2), .A1 (nx65890), .S0 (
             nx63550)) ;
    nand04 ix7823 (.Y (nx7822), .A0 (nx57634), .A1 (nx57642), .A2 (nx57650), .A3 (
           nx57658)) ;
    aoi22 ix57635 (.Y (nx57634), .A0 (ram_152__2), .A1 (nx64804), .B0 (
          ram_153__2), .B1 (nx64842)) ;
    dffr reg_ram_152__2 (.Q (ram_152__2), .QB (\$dummy [728]), .D (nx39140), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39141 (.Y (nx39140), .A0 (ram_152__2), .A1 (nx65890), .S0 (
             nx63542)) ;
    dffr reg_ram_153__2 (.Q (ram_153__2), .QB (\$dummy [729]), .D (nx39130), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39131 (.Y (nx39130), .A0 (ram_153__2), .A1 (nx65892), .S0 (
             nx63538)) ;
    aoi22 ix57643 (.Y (nx57642), .A0 (ram_155__2), .A1 (nx64880), .B0 (
          ram_154__2), .B1 (nx64918)) ;
    dffr reg_ram_155__2 (.Q (ram_155__2), .QB (\$dummy [730]), .D (nx39110), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39111 (.Y (nx39110), .A0 (ram_155__2), .A1 (nx65892), .S0 (
             nx63530)) ;
    dffr reg_ram_154__2 (.Q (ram_154__2), .QB (\$dummy [731]), .D (nx39120), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39121 (.Y (nx39120), .A0 (ram_154__2), .A1 (nx65892), .S0 (
             nx63534)) ;
    aoi22 ix57651 (.Y (nx57650), .A0 (ram_156__2), .A1 (nx64956), .B0 (
          ram_157__2), .B1 (nx64994)) ;
    dffr reg_ram_156__2 (.Q (ram_156__2), .QB (\$dummy [732]), .D (nx39100), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39101 (.Y (nx39100), .A0 (ram_156__2), .A1 (nx65892), .S0 (
             nx63526)) ;
    dffr reg_ram_157__2 (.Q (ram_157__2), .QB (\$dummy [733]), .D (nx39090), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39091 (.Y (nx39090), .A0 (ram_157__2), .A1 (nx65892), .S0 (
             nx63522)) ;
    aoi22 ix57659 (.Y (nx57658), .A0 (ram_159__2), .A1 (nx65032), .B0 (
          ram_158__2), .B1 (nx65070)) ;
    dffr reg_ram_159__2 (.Q (ram_159__2), .QB (\$dummy [734]), .D (nx39070), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39071 (.Y (nx39070), .A0 (ram_159__2), .A1 (nx65892), .S0 (
             nx63514)) ;
    dffr reg_ram_158__2 (.Q (ram_158__2), .QB (\$dummy [735]), .D (nx39080), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39081 (.Y (nx39080), .A0 (ram_158__2), .A1 (nx65892), .S0 (
             nx63518)) ;
    oai21 ix57667 (.Y (nx57666), .A0 (nx7736), .A1 (nx7658), .B0 (nx65222)) ;
    nand04 ix7737 (.Y (nx7736), .A0 (nx57669), .A1 (nx57677), .A2 (nx57685), .A3 (
           nx57693)) ;
    aoi22 ix57670 (.Y (nx57669), .A0 (ram_160__2), .A1 (nx64500), .B0 (
          ram_161__2), .B1 (nx64538)) ;
    dffr reg_ram_160__2 (.Q (ram_160__2), .QB (\$dummy [736]), .D (nx39060), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39061 (.Y (nx39060), .A0 (ram_160__2), .A1 (nx65894), .S0 (
             nx63504)) ;
    dffr reg_ram_161__2 (.Q (ram_161__2), .QB (\$dummy [737]), .D (nx39050), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39051 (.Y (nx39050), .A0 (ram_161__2), .A1 (nx65894), .S0 (
             nx63500)) ;
    aoi22 ix57678 (.Y (nx57677), .A0 (ram_163__2), .A1 (nx64576), .B0 (
          ram_162__2), .B1 (nx64614)) ;
    dffr reg_ram_163__2 (.Q (ram_163__2), .QB (\$dummy [738]), .D (nx39030), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39031 (.Y (nx39030), .A0 (ram_163__2), .A1 (nx65894), .S0 (
             nx63492)) ;
    dffr reg_ram_162__2 (.Q (ram_162__2), .QB (\$dummy [739]), .D (nx39040), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39041 (.Y (nx39040), .A0 (ram_162__2), .A1 (nx65894), .S0 (
             nx63496)) ;
    aoi22 ix57686 (.Y (nx57685), .A0 (ram_164__2), .A1 (nx64652), .B0 (
          ram_165__2), .B1 (nx64690)) ;
    dffr reg_ram_164__2 (.Q (ram_164__2), .QB (\$dummy [740]), .D (nx39020), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39021 (.Y (nx39020), .A0 (ram_164__2), .A1 (nx65894), .S0 (
             nx63488)) ;
    dffr reg_ram_165__2 (.Q (ram_165__2), .QB (\$dummy [741]), .D (nx39010), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39011 (.Y (nx39010), .A0 (ram_165__2), .A1 (nx65894), .S0 (
             nx63484)) ;
    aoi22 ix57694 (.Y (nx57693), .A0 (ram_167__2), .A1 (nx64728), .B0 (
          ram_166__2), .B1 (nx64766)) ;
    dffr reg_ram_167__2 (.Q (ram_167__2), .QB (\$dummy [742]), .D (nx38990), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38991 (.Y (nx38990), .A0 (ram_167__2), .A1 (nx65894), .S0 (
             nx63476)) ;
    dffr reg_ram_166__2 (.Q (ram_166__2), .QB (\$dummy [743]), .D (nx39000), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix39001 (.Y (nx39000), .A0 (ram_166__2), .A1 (nx65896), .S0 (
             nx63480)) ;
    nand04 ix7659 (.Y (nx7658), .A0 (nx57702), .A1 (nx57710), .A2 (nx57718), .A3 (
           nx57726)) ;
    aoi22 ix57703 (.Y (nx57702), .A0 (ram_168__2), .A1 (nx64804), .B0 (
          ram_169__2), .B1 (nx64842)) ;
    dffr reg_ram_168__2 (.Q (ram_168__2), .QB (\$dummy [744]), .D (nx38980), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38981 (.Y (nx38980), .A0 (ram_168__2), .A1 (nx65896), .S0 (
             nx63472)) ;
    dffr reg_ram_169__2 (.Q (ram_169__2), .QB (\$dummy [745]), .D (nx38970), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38971 (.Y (nx38970), .A0 (ram_169__2), .A1 (nx65896), .S0 (
             nx63468)) ;
    aoi22 ix57711 (.Y (nx57710), .A0 (ram_171__2), .A1 (nx64880), .B0 (
          ram_170__2), .B1 (nx64918)) ;
    dffr reg_ram_171__2 (.Q (ram_171__2), .QB (\$dummy [746]), .D (nx38950), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38951 (.Y (nx38950), .A0 (ram_171__2), .A1 (nx65896), .S0 (
             nx63460)) ;
    dffr reg_ram_170__2 (.Q (ram_170__2), .QB (\$dummy [747]), .D (nx38960), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38961 (.Y (nx38960), .A0 (ram_170__2), .A1 (nx65896), .S0 (
             nx63464)) ;
    aoi22 ix57719 (.Y (nx57718), .A0 (ram_172__2), .A1 (nx64956), .B0 (
          ram_173__2), .B1 (nx64994)) ;
    dffr reg_ram_172__2 (.Q (ram_172__2), .QB (\$dummy [748]), .D (nx38940), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38941 (.Y (nx38940), .A0 (ram_172__2), .A1 (nx65896), .S0 (
             nx63456)) ;
    dffr reg_ram_173__2 (.Q (ram_173__2), .QB (\$dummy [749]), .D (nx38930), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38931 (.Y (nx38930), .A0 (ram_173__2), .A1 (nx65896), .S0 (
             nx63452)) ;
    aoi22 ix57727 (.Y (nx57726), .A0 (ram_175__2), .A1 (nx65032), .B0 (
          ram_174__2), .B1 (nx65070)) ;
    dffr reg_ram_175__2 (.Q (ram_175__2), .QB (\$dummy [750]), .D (nx38910), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38911 (.Y (nx38910), .A0 (ram_175__2), .A1 (nx65898), .S0 (
             nx63444)) ;
    dffr reg_ram_174__2 (.Q (ram_174__2), .QB (\$dummy [751]), .D (nx38920), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38921 (.Y (nx38920), .A0 (ram_174__2), .A1 (nx65898), .S0 (
             nx63448)) ;
    oai21 ix57735 (.Y (nx57734), .A0 (nx7574), .A1 (nx7496), .B0 (nx65226)) ;
    nand04 ix7575 (.Y (nx7574), .A0 (nx57737), .A1 (nx57745), .A2 (nx57753), .A3 (
           nx57761)) ;
    aoi22 ix57738 (.Y (nx57737), .A0 (ram_176__2), .A1 (nx64500), .B0 (
          ram_177__2), .B1 (nx64538)) ;
    dffr reg_ram_176__2 (.Q (ram_176__2), .QB (\$dummy [752]), .D (nx38900), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38901 (.Y (nx38900), .A0 (ram_176__2), .A1 (nx65898), .S0 (
             nx63434)) ;
    dffr reg_ram_177__2 (.Q (ram_177__2), .QB (\$dummy [753]), .D (nx38890), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38891 (.Y (nx38890), .A0 (ram_177__2), .A1 (nx65898), .S0 (
             nx63424)) ;
    aoi22 ix57746 (.Y (nx57745), .A0 (ram_179__2), .A1 (nx64576), .B0 (
          ram_178__2), .B1 (nx64614)) ;
    dffr reg_ram_179__2 (.Q (ram_179__2), .QB (\$dummy [754]), .D (nx38870), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38871 (.Y (nx38870), .A0 (ram_179__2), .A1 (nx65898), .S0 (
             nx63404)) ;
    dffr reg_ram_178__2 (.Q (ram_178__2), .QB (\$dummy [755]), .D (nx38880), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38881 (.Y (nx38880), .A0 (ram_178__2), .A1 (nx65898), .S0 (
             nx63414)) ;
    aoi22 ix57754 (.Y (nx57753), .A0 (ram_180__2), .A1 (nx64652), .B0 (
          ram_181__2), .B1 (nx64690)) ;
    dffr reg_ram_180__2 (.Q (ram_180__2), .QB (\$dummy [756]), .D (nx38860), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38861 (.Y (nx38860), .A0 (ram_180__2), .A1 (nx65898), .S0 (
             nx63394)) ;
    dffr reg_ram_181__2 (.Q (ram_181__2), .QB (\$dummy [757]), .D (nx38850), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38851 (.Y (nx38850), .A0 (ram_181__2), .A1 (nx65900), .S0 (
             nx63384)) ;
    aoi22 ix57762 (.Y (nx57761), .A0 (ram_183__2), .A1 (nx64728), .B0 (
          ram_182__2), .B1 (nx64766)) ;
    dffr reg_ram_183__2 (.Q (ram_183__2), .QB (\$dummy [758]), .D (nx38830), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38831 (.Y (nx38830), .A0 (ram_183__2), .A1 (nx65900), .S0 (
             nx63364)) ;
    dffr reg_ram_182__2 (.Q (ram_182__2), .QB (\$dummy [759]), .D (nx38840), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38841 (.Y (nx38840), .A0 (ram_182__2), .A1 (nx65900), .S0 (
             nx63374)) ;
    nand04 ix7497 (.Y (nx7496), .A0 (nx57770), .A1 (nx57778), .A2 (nx57786), .A3 (
           nx57794)) ;
    aoi22 ix57771 (.Y (nx57770), .A0 (ram_184__2), .A1 (nx64804), .B0 (
          ram_185__2), .B1 (nx64842)) ;
    dffr reg_ram_184__2 (.Q (ram_184__2), .QB (\$dummy [760]), .D (nx38820), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38821 (.Y (nx38820), .A0 (ram_184__2), .A1 (nx65900), .S0 (
             nx63354)) ;
    dffr reg_ram_185__2 (.Q (ram_185__2), .QB (\$dummy [761]), .D (nx38810), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38811 (.Y (nx38810), .A0 (ram_185__2), .A1 (nx65900), .S0 (
             nx63344)) ;
    aoi22 ix57779 (.Y (nx57778), .A0 (ram_187__2), .A1 (nx64880), .B0 (
          ram_186__2), .B1 (nx64918)) ;
    dffr reg_ram_187__2 (.Q (ram_187__2), .QB (\$dummy [762]), .D (nx38790), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38791 (.Y (nx38790), .A0 (ram_187__2), .A1 (nx65900), .S0 (
             nx63324)) ;
    dffr reg_ram_186__2 (.Q (ram_186__2), .QB (\$dummy [763]), .D (nx38800), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38801 (.Y (nx38800), .A0 (ram_186__2), .A1 (nx65900), .S0 (
             nx63334)) ;
    aoi22 ix57787 (.Y (nx57786), .A0 (ram_188__2), .A1 (nx64956), .B0 (
          ram_189__2), .B1 (nx64994)) ;
    dffr reg_ram_188__2 (.Q (ram_188__2), .QB (\$dummy [764]), .D (nx38780), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38781 (.Y (nx38780), .A0 (ram_188__2), .A1 (nx65902), .S0 (
             nx63314)) ;
    dffr reg_ram_189__2 (.Q (ram_189__2), .QB (\$dummy [765]), .D (nx38770), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38771 (.Y (nx38770), .A0 (ram_189__2), .A1 (nx65902), .S0 (
             nx63304)) ;
    aoi22 ix57795 (.Y (nx57794), .A0 (ram_191__2), .A1 (nx65032), .B0 (
          ram_190__2), .B1 (nx65070)) ;
    dffr reg_ram_191__2 (.Q (ram_191__2), .QB (\$dummy [766]), .D (nx38750), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38751 (.Y (nx38750), .A0 (ram_191__2), .A1 (nx65902), .S0 (
             nx63284)) ;
    dffr reg_ram_190__2 (.Q (ram_190__2), .QB (\$dummy [767]), .D (nx38760), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix38761 (.Y (nx38760), .A0 (ram_190__2), .A1 (nx65902), .S0 (
             nx63294)) ;
    or04 ix12663 (.Y (dataout[3]), .A0 (nx12658), .A1 (nx12004), .A2 (nx11348), 
         .A3 (nx10694)) ;
    nand04 ix12659 (.Y (nx12658), .A0 (nx57804), .A1 (nx57872), .A2 (nx57940), .A3 (
           nx58008)) ;
    oai21 ix57805 (.Y (nx57804), .A0 (nx12648), .A1 (nx12570), .B0 (nx65096)) ;
    nand04 ix12649 (.Y (nx12648), .A0 (nx57807), .A1 (nx57815), .A2 (nx57823), .A3 (
           nx57831)) ;
    aoi22 ix57808 (.Y (nx57807), .A0 (ram_240__3), .A1 (nx64502), .B0 (
          ram_241__3), .B1 (nx64540)) ;
    dffr reg_ram_240__3 (.Q (ram_240__3), .QB (\$dummy [768]), .D (nx43860), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43861 (.Y (nx43860), .A0 (ram_240__3), .A1 (nx65754), .S0 (
             nx64414)) ;
    dffr reg_ram_241__3 (.Q (ram_241__3), .QB (\$dummy [769]), .D (nx43850), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43851 (.Y (nx43850), .A0 (ram_241__3), .A1 (nx65754), .S0 (
             nx64410)) ;
    aoi22 ix57816 (.Y (nx57815), .A0 (ram_243__3), .A1 (nx64578), .B0 (
          ram_242__3), .B1 (nx64616)) ;
    dffr reg_ram_243__3 (.Q (ram_243__3), .QB (\$dummy [770]), .D (nx43830), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43831 (.Y (nx43830), .A0 (ram_243__3), .A1 (nx65754), .S0 (
             nx64402)) ;
    dffr reg_ram_242__3 (.Q (ram_242__3), .QB (\$dummy [771]), .D (nx43840), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43841 (.Y (nx43840), .A0 (ram_242__3), .A1 (nx65754), .S0 (
             nx64406)) ;
    aoi22 ix57824 (.Y (nx57823), .A0 (ram_244__3), .A1 (nx64654), .B0 (
          ram_245__3), .B1 (nx64692)) ;
    dffr reg_ram_244__3 (.Q (ram_244__3), .QB (\$dummy [772]), .D (nx43820), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43821 (.Y (nx43820), .A0 (ram_244__3), .A1 (nx65754), .S0 (
             nx64398)) ;
    dffr reg_ram_245__3 (.Q (ram_245__3), .QB (\$dummy [773]), .D (nx43810), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43811 (.Y (nx43810), .A0 (ram_245__3), .A1 (nx65754), .S0 (
             nx64394)) ;
    aoi22 ix57832 (.Y (nx57831), .A0 (ram_247__3), .A1 (nx64730), .B0 (
          ram_246__3), .B1 (nx64768)) ;
    dffr reg_ram_247__3 (.Q (ram_247__3), .QB (\$dummy [774]), .D (nx43790), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43791 (.Y (nx43790), .A0 (ram_247__3), .A1 (nx65754), .S0 (
             nx64386)) ;
    dffr reg_ram_246__3 (.Q (ram_246__3), .QB (\$dummy [775]), .D (nx43800), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43801 (.Y (nx43800), .A0 (ram_246__3), .A1 (nx65756), .S0 (
             nx64390)) ;
    nand04 ix12571 (.Y (nx12570), .A0 (nx57840), .A1 (nx57848), .A2 (nx57856), .A3 (
           nx57864)) ;
    aoi22 ix57841 (.Y (nx57840), .A0 (ram_248__3), .A1 (nx64806), .B0 (
          ram_249__3), .B1 (nx64844)) ;
    dffr reg_ram_248__3 (.Q (ram_248__3), .QB (\$dummy [776]), .D (nx43780), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43781 (.Y (nx43780), .A0 (ram_248__3), .A1 (nx65756), .S0 (
             nx64382)) ;
    dffr reg_ram_249__3 (.Q (ram_249__3), .QB (\$dummy [777]), .D (nx43770), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43771 (.Y (nx43770), .A0 (ram_249__3), .A1 (nx65756), .S0 (
             nx64378)) ;
    aoi22 ix57849 (.Y (nx57848), .A0 (ram_251__3), .A1 (nx64882), .B0 (
          ram_250__3), .B1 (nx64920)) ;
    dffr reg_ram_251__3 (.Q (ram_251__3), .QB (\$dummy [778]), .D (nx43750), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43751 (.Y (nx43750), .A0 (ram_251__3), .A1 (nx65756), .S0 (
             nx64370)) ;
    dffr reg_ram_250__3 (.Q (ram_250__3), .QB (\$dummy [779]), .D (nx43760), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43761 (.Y (nx43760), .A0 (ram_250__3), .A1 (nx65756), .S0 (
             nx64374)) ;
    aoi22 ix57857 (.Y (nx57856), .A0 (ram_252__3), .A1 (nx64958), .B0 (
          ram_253__3), .B1 (nx64996)) ;
    dffr reg_ram_252__3 (.Q (ram_252__3), .QB (\$dummy [780]), .D (nx43740), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43741 (.Y (nx43740), .A0 (ram_252__3), .A1 (nx65756), .S0 (
             nx64366)) ;
    dffr reg_ram_253__3 (.Q (ram_253__3), .QB (\$dummy [781]), .D (nx43730), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43731 (.Y (nx43730), .A0 (ram_253__3), .A1 (nx65756), .S0 (
             nx64362)) ;
    aoi22 ix57865 (.Y (nx57864), .A0 (ram_255__3), .A1 (nx65034), .B0 (
          ram_254__3), .B1 (nx65072)) ;
    dffr reg_ram_255__3 (.Q (ram_255__3), .QB (\$dummy [782]), .D (nx43710), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43711 (.Y (nx43710), .A0 (ram_255__3), .A1 (nx65758), .S0 (
             nx64354)) ;
    dffr reg_ram_254__3 (.Q (ram_254__3), .QB (\$dummy [783]), .D (nx43720), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43721 (.Y (nx43720), .A0 (ram_254__3), .A1 (nx65758), .S0 (
             nx64358)) ;
    oai21 ix57873 (.Y (nx57872), .A0 (nx12486), .A1 (nx12408), .B0 (nx65100)) ;
    nand04 ix12487 (.Y (nx12486), .A0 (nx57875), .A1 (nx57883), .A2 (nx57891), .A3 (
           nx57899)) ;
    aoi22 ix57876 (.Y (nx57875), .A0 (ram_224__3), .A1 (nx64502), .B0 (
          ram_225__3), .B1 (nx64540)) ;
    dffr reg_ram_224__3 (.Q (ram_224__3), .QB (\$dummy [784]), .D (nx43700), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43701 (.Y (nx43700), .A0 (ram_224__3), .A1 (nx65758), .S0 (
             nx64344)) ;
    dffr reg_ram_225__3 (.Q (ram_225__3), .QB (\$dummy [785]), .D (nx43690), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43691 (.Y (nx43690), .A0 (ram_225__3), .A1 (nx65758), .S0 (
             nx64340)) ;
    aoi22 ix57884 (.Y (nx57883), .A0 (ram_227__3), .A1 (nx64578), .B0 (
          ram_226__3), .B1 (nx64616)) ;
    dffr reg_ram_227__3 (.Q (ram_227__3), .QB (\$dummy [786]), .D (nx43670), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43671 (.Y (nx43670), .A0 (ram_227__3), .A1 (nx65758), .S0 (
             nx64332)) ;
    dffr reg_ram_226__3 (.Q (ram_226__3), .QB (\$dummy [787]), .D (nx43680), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43681 (.Y (nx43680), .A0 (ram_226__3), .A1 (nx65758), .S0 (
             nx64336)) ;
    aoi22 ix57892 (.Y (nx57891), .A0 (ram_228__3), .A1 (nx64654), .B0 (
          ram_229__3), .B1 (nx64692)) ;
    dffr reg_ram_228__3 (.Q (ram_228__3), .QB (\$dummy [788]), .D (nx43660), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43661 (.Y (nx43660), .A0 (ram_228__3), .A1 (nx65758), .S0 (
             nx64328)) ;
    dffr reg_ram_229__3 (.Q (ram_229__3), .QB (\$dummy [789]), .D (nx43650), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43651 (.Y (nx43650), .A0 (ram_229__3), .A1 (nx65760), .S0 (
             nx64324)) ;
    aoi22 ix57900 (.Y (nx57899), .A0 (ram_231__3), .A1 (nx64730), .B0 (
          ram_230__3), .B1 (nx64768)) ;
    dffr reg_ram_231__3 (.Q (ram_231__3), .QB (\$dummy [790]), .D (nx43630), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43631 (.Y (nx43630), .A0 (ram_231__3), .A1 (nx65760), .S0 (
             nx64316)) ;
    dffr reg_ram_230__3 (.Q (ram_230__3), .QB (\$dummy [791]), .D (nx43640), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43641 (.Y (nx43640), .A0 (ram_230__3), .A1 (nx65760), .S0 (
             nx64320)) ;
    nand04 ix12409 (.Y (nx12408), .A0 (nx57908), .A1 (nx57916), .A2 (nx57924), .A3 (
           nx57932)) ;
    aoi22 ix57909 (.Y (nx57908), .A0 (ram_232__3), .A1 (nx64806), .B0 (
          ram_233__3), .B1 (nx64844)) ;
    dffr reg_ram_232__3 (.Q (ram_232__3), .QB (\$dummy [792]), .D (nx43620), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43621 (.Y (nx43620), .A0 (ram_232__3), .A1 (nx65760), .S0 (
             nx64312)) ;
    dffr reg_ram_233__3 (.Q (ram_233__3), .QB (\$dummy [793]), .D (nx43610), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43611 (.Y (nx43610), .A0 (ram_233__3), .A1 (nx65760), .S0 (
             nx64308)) ;
    aoi22 ix57917 (.Y (nx57916), .A0 (ram_235__3), .A1 (nx64882), .B0 (
          ram_234__3), .B1 (nx64920)) ;
    dffr reg_ram_235__3 (.Q (ram_235__3), .QB (\$dummy [794]), .D (nx43590), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43591 (.Y (nx43590), .A0 (ram_235__3), .A1 (nx65760), .S0 (
             nx64300)) ;
    dffr reg_ram_234__3 (.Q (ram_234__3), .QB (\$dummy [795]), .D (nx43600), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43601 (.Y (nx43600), .A0 (ram_234__3), .A1 (nx65760), .S0 (
             nx64304)) ;
    aoi22 ix57925 (.Y (nx57924), .A0 (ram_236__3), .A1 (nx64958), .B0 (
          ram_237__3), .B1 (nx64996)) ;
    dffr reg_ram_236__3 (.Q (ram_236__3), .QB (\$dummy [796]), .D (nx43580), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43581 (.Y (nx43580), .A0 (ram_236__3), .A1 (nx65762), .S0 (
             nx64296)) ;
    dffr reg_ram_237__3 (.Q (ram_237__3), .QB (\$dummy [797]), .D (nx43570), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43571 (.Y (nx43570), .A0 (ram_237__3), .A1 (nx65762), .S0 (
             nx64292)) ;
    aoi22 ix57933 (.Y (nx57932), .A0 (ram_239__3), .A1 (nx65034), .B0 (
          ram_238__3), .B1 (nx65072)) ;
    dffr reg_ram_239__3 (.Q (ram_239__3), .QB (\$dummy [798]), .D (nx43550), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43551 (.Y (nx43550), .A0 (ram_239__3), .A1 (nx65762), .S0 (
             nx64284)) ;
    dffr reg_ram_238__3 (.Q (ram_238__3), .QB (\$dummy [799]), .D (nx43560), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43561 (.Y (nx43560), .A0 (ram_238__3), .A1 (nx65762), .S0 (
             nx64288)) ;
    oai21 ix57941 (.Y (nx57940), .A0 (nx12322), .A1 (nx12244), .B0 (nx65104)) ;
    nand04 ix12323 (.Y (nx12322), .A0 (nx57943), .A1 (nx57951), .A2 (nx57959), .A3 (
           nx57967)) ;
    aoi22 ix57944 (.Y (nx57943), .A0 (ram_208__3), .A1 (nx64502), .B0 (
          ram_209__3), .B1 (nx64540)) ;
    dffr reg_ram_208__3 (.Q (ram_208__3), .QB (\$dummy [800]), .D (nx43540), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43541 (.Y (nx43540), .A0 (ram_208__3), .A1 (nx65762), .S0 (
             nx64274)) ;
    dffr reg_ram_209__3 (.Q (ram_209__3), .QB (\$dummy [801]), .D (nx43530), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43531 (.Y (nx43530), .A0 (ram_209__3), .A1 (nx65762), .S0 (
             nx64270)) ;
    aoi22 ix57952 (.Y (nx57951), .A0 (ram_211__3), .A1 (nx64578), .B0 (
          ram_210__3), .B1 (nx64616)) ;
    dffr reg_ram_211__3 (.Q (ram_211__3), .QB (\$dummy [802]), .D (nx43510), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43511 (.Y (nx43510), .A0 (ram_211__3), .A1 (nx65762), .S0 (
             nx64262)) ;
    dffr reg_ram_210__3 (.Q (ram_210__3), .QB (\$dummy [803]), .D (nx43520), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43521 (.Y (nx43520), .A0 (ram_210__3), .A1 (nx65764), .S0 (
             nx64266)) ;
    aoi22 ix57960 (.Y (nx57959), .A0 (ram_212__3), .A1 (nx64654), .B0 (
          ram_213__3), .B1 (nx64692)) ;
    dffr reg_ram_212__3 (.Q (ram_212__3), .QB (\$dummy [804]), .D (nx43500), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43501 (.Y (nx43500), .A0 (ram_212__3), .A1 (nx65764), .S0 (
             nx64258)) ;
    dffr reg_ram_213__3 (.Q (ram_213__3), .QB (\$dummy [805]), .D (nx43490), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43491 (.Y (nx43490), .A0 (ram_213__3), .A1 (nx65764), .S0 (
             nx64254)) ;
    aoi22 ix57968 (.Y (nx57967), .A0 (ram_215__3), .A1 (nx64730), .B0 (
          ram_214__3), .B1 (nx64768)) ;
    dffr reg_ram_215__3 (.Q (ram_215__3), .QB (\$dummy [806]), .D (nx43470), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43471 (.Y (nx43470), .A0 (ram_215__3), .A1 (nx65764), .S0 (
             nx64246)) ;
    dffr reg_ram_214__3 (.Q (ram_214__3), .QB (\$dummy [807]), .D (nx43480), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43481 (.Y (nx43480), .A0 (ram_214__3), .A1 (nx65764), .S0 (
             nx64250)) ;
    nand04 ix12245 (.Y (nx12244), .A0 (nx57976), .A1 (nx57984), .A2 (nx57992), .A3 (
           nx58000)) ;
    aoi22 ix57977 (.Y (nx57976), .A0 (ram_216__3), .A1 (nx64806), .B0 (
          ram_217__3), .B1 (nx64844)) ;
    dffr reg_ram_216__3 (.Q (ram_216__3), .QB (\$dummy [808]), .D (nx43460), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43461 (.Y (nx43460), .A0 (ram_216__3), .A1 (nx65764), .S0 (
             nx64242)) ;
    dffr reg_ram_217__3 (.Q (ram_217__3), .QB (\$dummy [809]), .D (nx43450), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43451 (.Y (nx43450), .A0 (ram_217__3), .A1 (nx65764), .S0 (
             nx64238)) ;
    aoi22 ix57985 (.Y (nx57984), .A0 (ram_219__3), .A1 (nx64882), .B0 (
          ram_218__3), .B1 (nx64920)) ;
    dffr reg_ram_219__3 (.Q (ram_219__3), .QB (\$dummy [810]), .D (nx43430), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43431 (.Y (nx43430), .A0 (ram_219__3), .A1 (nx65766), .S0 (
             nx64230)) ;
    dffr reg_ram_218__3 (.Q (ram_218__3), .QB (\$dummy [811]), .D (nx43440), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43441 (.Y (nx43440), .A0 (ram_218__3), .A1 (nx65766), .S0 (
             nx64234)) ;
    aoi22 ix57993 (.Y (nx57992), .A0 (ram_220__3), .A1 (nx64958), .B0 (
          ram_221__3), .B1 (nx64996)) ;
    dffr reg_ram_220__3 (.Q (ram_220__3), .QB (\$dummy [812]), .D (nx43420), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43421 (.Y (nx43420), .A0 (ram_220__3), .A1 (nx65766), .S0 (
             nx64226)) ;
    dffr reg_ram_221__3 (.Q (ram_221__3), .QB (\$dummy [813]), .D (nx43410), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43411 (.Y (nx43410), .A0 (ram_221__3), .A1 (nx65766), .S0 (
             nx64222)) ;
    aoi22 ix58001 (.Y (nx58000), .A0 (ram_223__3), .A1 (nx65034), .B0 (
          ram_222__3), .B1 (nx65072)) ;
    dffr reg_ram_223__3 (.Q (ram_223__3), .QB (\$dummy [814]), .D (nx43390), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43391 (.Y (nx43390), .A0 (ram_223__3), .A1 (nx65766), .S0 (
             nx64214)) ;
    dffr reg_ram_222__3 (.Q (ram_222__3), .QB (\$dummy [815]), .D (nx43400), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43401 (.Y (nx43400), .A0 (ram_222__3), .A1 (nx65766), .S0 (
             nx64218)) ;
    oai21 ix58009 (.Y (nx58008), .A0 (nx12160), .A1 (nx12082), .B0 (nx65108)) ;
    nand04 ix12161 (.Y (nx12160), .A0 (nx58011), .A1 (nx58019), .A2 (nx58027), .A3 (
           nx58035)) ;
    aoi22 ix58012 (.Y (nx58011), .A0 (ram_192__3), .A1 (nx64502), .B0 (
          ram_193__3), .B1 (nx64540)) ;
    dffr reg_ram_192__3 (.Q (ram_192__3), .QB (\$dummy [816]), .D (nx43380), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43381 (.Y (nx43380), .A0 (ram_192__3), .A1 (nx65766), .S0 (
             nx64204)) ;
    dffr reg_ram_193__3 (.Q (ram_193__3), .QB (\$dummy [817]), .D (nx43370), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43371 (.Y (nx43370), .A0 (ram_193__3), .A1 (nx65768), .S0 (
             nx64200)) ;
    aoi22 ix58020 (.Y (nx58019), .A0 (ram_195__3), .A1 (nx64578), .B0 (
          ram_194__3), .B1 (nx64616)) ;
    dffr reg_ram_195__3 (.Q (ram_195__3), .QB (\$dummy [818]), .D (nx43350), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43351 (.Y (nx43350), .A0 (ram_195__3), .A1 (nx65768), .S0 (
             nx64192)) ;
    dffr reg_ram_194__3 (.Q (ram_194__3), .QB (\$dummy [819]), .D (nx43360), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43361 (.Y (nx43360), .A0 (ram_194__3), .A1 (nx65768), .S0 (
             nx64196)) ;
    aoi22 ix58028 (.Y (nx58027), .A0 (ram_196__3), .A1 (nx64654), .B0 (
          ram_197__3), .B1 (nx64692)) ;
    dffr reg_ram_196__3 (.Q (ram_196__3), .QB (\$dummy [820]), .D (nx43340), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43341 (.Y (nx43340), .A0 (ram_196__3), .A1 (nx65768), .S0 (
             nx64188)) ;
    dffr reg_ram_197__3 (.Q (ram_197__3), .QB (\$dummy [821]), .D (nx43330), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43331 (.Y (nx43330), .A0 (ram_197__3), .A1 (nx65768), .S0 (
             nx64184)) ;
    aoi22 ix58036 (.Y (nx58035), .A0 (ram_199__3), .A1 (nx64730), .B0 (
          ram_198__3), .B1 (nx64768)) ;
    dffr reg_ram_199__3 (.Q (ram_199__3), .QB (\$dummy [822]), .D (nx43310), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43311 (.Y (nx43310), .A0 (ram_199__3), .A1 (nx65768), .S0 (
             nx64176)) ;
    dffr reg_ram_198__3 (.Q (ram_198__3), .QB (\$dummy [823]), .D (nx43320), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43321 (.Y (nx43320), .A0 (ram_198__3), .A1 (nx65768), .S0 (
             nx64180)) ;
    nand04 ix12083 (.Y (nx12082), .A0 (nx58044), .A1 (nx58052), .A2 (nx58060), .A3 (
           nx58068)) ;
    aoi22 ix58045 (.Y (nx58044), .A0 (ram_200__3), .A1 (nx64806), .B0 (
          ram_201__3), .B1 (nx64844)) ;
    dffr reg_ram_200__3 (.Q (ram_200__3), .QB (\$dummy [824]), .D (nx43300), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43301 (.Y (nx43300), .A0 (ram_200__3), .A1 (nx65770), .S0 (
             nx64172)) ;
    dffr reg_ram_201__3 (.Q (ram_201__3), .QB (\$dummy [825]), .D (nx43290), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43291 (.Y (nx43290), .A0 (ram_201__3), .A1 (nx65770), .S0 (
             nx64168)) ;
    aoi22 ix58053 (.Y (nx58052), .A0 (ram_203__3), .A1 (nx64882), .B0 (
          ram_202__3), .B1 (nx64920)) ;
    dffr reg_ram_203__3 (.Q (ram_203__3), .QB (\$dummy [826]), .D (nx43270), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43271 (.Y (nx43270), .A0 (ram_203__3), .A1 (nx65770), .S0 (
             nx64160)) ;
    dffr reg_ram_202__3 (.Q (ram_202__3), .QB (\$dummy [827]), .D (nx43280), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43281 (.Y (nx43280), .A0 (ram_202__3), .A1 (nx65770), .S0 (
             nx64164)) ;
    aoi22 ix58061 (.Y (nx58060), .A0 (ram_204__3), .A1 (nx64958), .B0 (
          ram_205__3), .B1 (nx64996)) ;
    dffr reg_ram_204__3 (.Q (ram_204__3), .QB (\$dummy [828]), .D (nx43260), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43261 (.Y (nx43260), .A0 (ram_204__3), .A1 (nx65770), .S0 (
             nx64156)) ;
    dffr reg_ram_205__3 (.Q (ram_205__3), .QB (\$dummy [829]), .D (nx43250), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43251 (.Y (nx43250), .A0 (ram_205__3), .A1 (nx65770), .S0 (
             nx64152)) ;
    aoi22 ix58069 (.Y (nx58068), .A0 (ram_207__3), .A1 (nx65034), .B0 (
          ram_206__3), .B1 (nx65072)) ;
    dffr reg_ram_207__3 (.Q (ram_207__3), .QB (\$dummy [830]), .D (nx43230), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43231 (.Y (nx43230), .A0 (ram_207__3), .A1 (nx65770), .S0 (
             nx64144)) ;
    dffr reg_ram_206__3 (.Q (ram_206__3), .QB (\$dummy [831]), .D (nx43240), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43241 (.Y (nx43240), .A0 (ram_206__3), .A1 (nx65772), .S0 (
             nx64148)) ;
    nand04 ix12005 (.Y (nx12004), .A0 (nx58077), .A1 (nx58145), .A2 (nx58213), .A3 (
           nx58281)) ;
    oai21 ix58078 (.Y (nx58077), .A0 (nx11994), .A1 (nx11916), .B0 (nx65112)) ;
    nand04 ix11995 (.Y (nx11994), .A0 (nx58080), .A1 (nx58088), .A2 (nx58096), .A3 (
           nx58104)) ;
    aoi22 ix58081 (.Y (nx58080), .A0 (ram_80__3), .A1 (nx64502), .B0 (ram_81__3)
          , .B1 (nx64540)) ;
    dffr reg_ram_80__3 (.Q (ram_80__3), .QB (\$dummy [832]), .D (nx43220), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43221 (.Y (nx43220), .A0 (ram_80__3), .A1 (nx65772), .S0 (nx64134
             )) ;
    dffr reg_ram_81__3 (.Q (ram_81__3), .QB (\$dummy [833]), .D (nx43210), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43211 (.Y (nx43210), .A0 (ram_81__3), .A1 (nx65772), .S0 (nx64130
             )) ;
    aoi22 ix58089 (.Y (nx58088), .A0 (ram_83__3), .A1 (nx64578), .B0 (ram_82__3)
          , .B1 (nx64616)) ;
    dffr reg_ram_83__3 (.Q (ram_83__3), .QB (\$dummy [834]), .D (nx43190), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43191 (.Y (nx43190), .A0 (ram_83__3), .A1 (nx65772), .S0 (nx64122
             )) ;
    dffr reg_ram_82__3 (.Q (ram_82__3), .QB (\$dummy [835]), .D (nx43200), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43201 (.Y (nx43200), .A0 (ram_82__3), .A1 (nx65772), .S0 (nx64126
             )) ;
    aoi22 ix58097 (.Y (nx58096), .A0 (ram_84__3), .A1 (nx64654), .B0 (ram_85__3)
          , .B1 (nx64692)) ;
    dffr reg_ram_84__3 (.Q (ram_84__3), .QB (\$dummy [836]), .D (nx43180), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43181 (.Y (nx43180), .A0 (ram_84__3), .A1 (nx65772), .S0 (nx64118
             )) ;
    dffr reg_ram_85__3 (.Q (ram_85__3), .QB (\$dummy [837]), .D (nx43170), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43171 (.Y (nx43170), .A0 (ram_85__3), .A1 (nx65772), .S0 (nx64114
             )) ;
    aoi22 ix58105 (.Y (nx58104), .A0 (ram_87__3), .A1 (nx64730), .B0 (ram_86__3)
          , .B1 (nx64768)) ;
    dffr reg_ram_87__3 (.Q (ram_87__3), .QB (\$dummy [838]), .D (nx43150), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43151 (.Y (nx43150), .A0 (ram_87__3), .A1 (nx65774), .S0 (nx64106
             )) ;
    dffr reg_ram_86__3 (.Q (ram_86__3), .QB (\$dummy [839]), .D (nx43160), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43161 (.Y (nx43160), .A0 (ram_86__3), .A1 (nx65774), .S0 (nx64110
             )) ;
    nand04 ix11917 (.Y (nx11916), .A0 (nx58113), .A1 (nx58121), .A2 (nx58129), .A3 (
           nx58137)) ;
    aoi22 ix58114 (.Y (nx58113), .A0 (ram_88__3), .A1 (nx64806), .B0 (ram_89__3)
          , .B1 (nx64844)) ;
    dffr reg_ram_88__3 (.Q (ram_88__3), .QB (\$dummy [840]), .D (nx43140), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43141 (.Y (nx43140), .A0 (ram_88__3), .A1 (nx65774), .S0 (nx64102
             )) ;
    dffr reg_ram_89__3 (.Q (ram_89__3), .QB (\$dummy [841]), .D (nx43130), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43131 (.Y (nx43130), .A0 (ram_89__3), .A1 (nx65774), .S0 (nx64098
             )) ;
    aoi22 ix58122 (.Y (nx58121), .A0 (ram_91__3), .A1 (nx64882), .B0 (ram_90__3)
          , .B1 (nx64920)) ;
    dffr reg_ram_91__3 (.Q (ram_91__3), .QB (\$dummy [842]), .D (nx43110), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43111 (.Y (nx43110), .A0 (ram_91__3), .A1 (nx65774), .S0 (nx64090
             )) ;
    dffr reg_ram_90__3 (.Q (ram_90__3), .QB (\$dummy [843]), .D (nx43120), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43121 (.Y (nx43120), .A0 (ram_90__3), .A1 (nx65774), .S0 (nx64094
             )) ;
    aoi22 ix58130 (.Y (nx58129), .A0 (ram_92__3), .A1 (nx64958), .B0 (ram_93__3)
          , .B1 (nx64996)) ;
    dffr reg_ram_92__3 (.Q (ram_92__3), .QB (\$dummy [844]), .D (nx43100), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43101 (.Y (nx43100), .A0 (ram_92__3), .A1 (nx65774), .S0 (nx64086
             )) ;
    dffr reg_ram_93__3 (.Q (ram_93__3), .QB (\$dummy [845]), .D (nx43090), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43091 (.Y (nx43090), .A0 (ram_93__3), .A1 (nx65776), .S0 (nx64082
             )) ;
    aoi22 ix58138 (.Y (nx58137), .A0 (ram_95__3), .A1 (nx65034), .B0 (ram_94__3)
          , .B1 (nx65072)) ;
    dffr reg_ram_95__3 (.Q (ram_95__3), .QB (\$dummy [846]), .D (nx43070), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43071 (.Y (nx43070), .A0 (ram_95__3), .A1 (nx65776), .S0 (nx64074
             )) ;
    dffr reg_ram_94__3 (.Q (ram_94__3), .QB (\$dummy [847]), .D (nx43080), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43081 (.Y (nx43080), .A0 (ram_94__3), .A1 (nx65776), .S0 (nx64078
             )) ;
    oai21 ix58146 (.Y (nx58145), .A0 (nx11832), .A1 (nx11754), .B0 (nx65116)) ;
    nand04 ix11833 (.Y (nx11832), .A0 (nx58148), .A1 (nx58156), .A2 (nx58164), .A3 (
           nx58172)) ;
    aoi22 ix58149 (.Y (nx58148), .A0 (ram_64__3), .A1 (nx64502), .B0 (ram_65__3)
          , .B1 (nx64540)) ;
    dffr reg_ram_64__3 (.Q (ram_64__3), .QB (\$dummy [848]), .D (nx43060), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43061 (.Y (nx43060), .A0 (ram_64__3), .A1 (nx65776), .S0 (nx64064
             )) ;
    dffr reg_ram_65__3 (.Q (ram_65__3), .QB (\$dummy [849]), .D (nx43050), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43051 (.Y (nx43050), .A0 (ram_65__3), .A1 (nx65776), .S0 (nx64060
             )) ;
    aoi22 ix58157 (.Y (nx58156), .A0 (ram_67__3), .A1 (nx64578), .B0 (ram_66__3)
          , .B1 (nx64616)) ;
    dffr reg_ram_67__3 (.Q (ram_67__3), .QB (\$dummy [850]), .D (nx43030), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43031 (.Y (nx43030), .A0 (ram_67__3), .A1 (nx65776), .S0 (nx64052
             )) ;
    dffr reg_ram_66__3 (.Q (ram_66__3), .QB (\$dummy [851]), .D (nx43040), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43041 (.Y (nx43040), .A0 (ram_66__3), .A1 (nx65776), .S0 (nx64056
             )) ;
    aoi22 ix58165 (.Y (nx58164), .A0 (ram_68__3), .A1 (nx64654), .B0 (ram_69__3)
          , .B1 (nx64692)) ;
    dffr reg_ram_68__3 (.Q (ram_68__3), .QB (\$dummy [852]), .D (nx43020), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43021 (.Y (nx43020), .A0 (ram_68__3), .A1 (nx65778), .S0 (nx64048
             )) ;
    dffr reg_ram_69__3 (.Q (ram_69__3), .QB (\$dummy [853]), .D (nx43010), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43011 (.Y (nx43010), .A0 (ram_69__3), .A1 (nx65778), .S0 (nx64044
             )) ;
    aoi22 ix58173 (.Y (nx58172), .A0 (ram_71__3), .A1 (nx64730), .B0 (ram_70__3)
          , .B1 (nx64768)) ;
    dffr reg_ram_71__3 (.Q (ram_71__3), .QB (\$dummy [854]), .D (nx42990), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42991 (.Y (nx42990), .A0 (ram_71__3), .A1 (nx65778), .S0 (nx64036
             )) ;
    dffr reg_ram_70__3 (.Q (ram_70__3), .QB (\$dummy [855]), .D (nx43000), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43001 (.Y (nx43000), .A0 (ram_70__3), .A1 (nx65778), .S0 (nx64040
             )) ;
    nand04 ix11755 (.Y (nx11754), .A0 (nx58181), .A1 (nx58189), .A2 (nx58197), .A3 (
           nx58205)) ;
    aoi22 ix58182 (.Y (nx58181), .A0 (ram_72__3), .A1 (nx64806), .B0 (ram_73__3)
          , .B1 (nx64844)) ;
    dffr reg_ram_72__3 (.Q (ram_72__3), .QB (\$dummy [856]), .D (nx42980), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42981 (.Y (nx42980), .A0 (ram_72__3), .A1 (nx65778), .S0 (nx64032
             )) ;
    dffr reg_ram_73__3 (.Q (ram_73__3), .QB (\$dummy [857]), .D (nx42970), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42971 (.Y (nx42970), .A0 (ram_73__3), .A1 (nx65778), .S0 (nx64028
             )) ;
    aoi22 ix58190 (.Y (nx58189), .A0 (ram_75__3), .A1 (nx64882), .B0 (ram_74__3)
          , .B1 (nx64920)) ;
    dffr reg_ram_75__3 (.Q (ram_75__3), .QB (\$dummy [858]), .D (nx42950), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42951 (.Y (nx42950), .A0 (ram_75__3), .A1 (nx65778), .S0 (nx64020
             )) ;
    dffr reg_ram_74__3 (.Q (ram_74__3), .QB (\$dummy [859]), .D (nx42960), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42961 (.Y (nx42960), .A0 (ram_74__3), .A1 (nx65780), .S0 (nx64024
             )) ;
    aoi22 ix58198 (.Y (nx58197), .A0 (ram_76__3), .A1 (nx64958), .B0 (ram_77__3)
          , .B1 (nx64996)) ;
    dffr reg_ram_76__3 (.Q (ram_76__3), .QB (\$dummy [860]), .D (nx42940), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42941 (.Y (nx42940), .A0 (ram_76__3), .A1 (nx65780), .S0 (nx64016
             )) ;
    dffr reg_ram_77__3 (.Q (ram_77__3), .QB (\$dummy [861]), .D (nx42930), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42931 (.Y (nx42930), .A0 (ram_77__3), .A1 (nx65780), .S0 (nx64012
             )) ;
    aoi22 ix58206 (.Y (nx58205), .A0 (ram_79__3), .A1 (nx65034), .B0 (ram_78__3)
          , .B1 (nx65072)) ;
    dffr reg_ram_79__3 (.Q (ram_79__3), .QB (\$dummy [862]), .D (nx42910), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42911 (.Y (nx42910), .A0 (ram_79__3), .A1 (nx65780), .S0 (nx64004
             )) ;
    dffr reg_ram_78__3 (.Q (ram_78__3), .QB (\$dummy [863]), .D (nx42920), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42921 (.Y (nx42920), .A0 (ram_78__3), .A1 (nx65780), .S0 (nx64008
             )) ;
    oai21 ix58214 (.Y (nx58213), .A0 (nx11668), .A1 (nx11590), .B0 (nx65120)) ;
    nand04 ix11669 (.Y (nx11668), .A0 (nx58216), .A1 (nx58224), .A2 (nx58232), .A3 (
           nx58240)) ;
    aoi22 ix58217 (.Y (nx58216), .A0 (ram_48__3), .A1 (nx64502), .B0 (ram_49__3)
          , .B1 (nx64540)) ;
    dffr reg_ram_48__3 (.Q (ram_48__3), .QB (\$dummy [864]), .D (nx42900), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42901 (.Y (nx42900), .A0 (ram_48__3), .A1 (nx65780), .S0 (nx63994
             )) ;
    dffr reg_ram_49__3 (.Q (ram_49__3), .QB (\$dummy [865]), .D (nx42890), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42891 (.Y (nx42890), .A0 (ram_49__3), .A1 (nx65780), .S0 (nx63990
             )) ;
    aoi22 ix58225 (.Y (nx58224), .A0 (ram_51__3), .A1 (nx64578), .B0 (ram_50__3)
          , .B1 (nx64616)) ;
    dffr reg_ram_51__3 (.Q (ram_51__3), .QB (\$dummy [866]), .D (nx42870), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42871 (.Y (nx42870), .A0 (ram_51__3), .A1 (nx65782), .S0 (nx63982
             )) ;
    dffr reg_ram_50__3 (.Q (ram_50__3), .QB (\$dummy [867]), .D (nx42880), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42881 (.Y (nx42880), .A0 (ram_50__3), .A1 (nx65782), .S0 (nx63986
             )) ;
    aoi22 ix58233 (.Y (nx58232), .A0 (ram_52__3), .A1 (nx64654), .B0 (ram_53__3)
          , .B1 (nx64692)) ;
    dffr reg_ram_52__3 (.Q (ram_52__3), .QB (\$dummy [868]), .D (nx42860), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42861 (.Y (nx42860), .A0 (ram_52__3), .A1 (nx65782), .S0 (nx63978
             )) ;
    dffr reg_ram_53__3 (.Q (ram_53__3), .QB (\$dummy [869]), .D (nx42850), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42851 (.Y (nx42850), .A0 (ram_53__3), .A1 (nx65782), .S0 (nx63974
             )) ;
    aoi22 ix58241 (.Y (nx58240), .A0 (ram_55__3), .A1 (nx64730), .B0 (ram_54__3)
          , .B1 (nx64768)) ;
    dffr reg_ram_55__3 (.Q (ram_55__3), .QB (\$dummy [870]), .D (nx42830), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42831 (.Y (nx42830), .A0 (ram_55__3), .A1 (nx65782), .S0 (nx63966
             )) ;
    dffr reg_ram_54__3 (.Q (ram_54__3), .QB (\$dummy [871]), .D (nx42840), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42841 (.Y (nx42840), .A0 (ram_54__3), .A1 (nx65782), .S0 (nx63970
             )) ;
    nand04 ix11591 (.Y (nx11590), .A0 (nx58249), .A1 (nx58257), .A2 (nx58265), .A3 (
           nx58273)) ;
    aoi22 ix58250 (.Y (nx58249), .A0 (ram_56__3), .A1 (nx64806), .B0 (ram_57__3)
          , .B1 (nx64844)) ;
    dffr reg_ram_56__3 (.Q (ram_56__3), .QB (\$dummy [872]), .D (nx42820), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42821 (.Y (nx42820), .A0 (ram_56__3), .A1 (nx65782), .S0 (nx63962
             )) ;
    dffr reg_ram_57__3 (.Q (ram_57__3), .QB (\$dummy [873]), .D (nx42810), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42811 (.Y (nx42810), .A0 (ram_57__3), .A1 (nx65784), .S0 (nx63958
             )) ;
    aoi22 ix58258 (.Y (nx58257), .A0 (ram_59__3), .A1 (nx64882), .B0 (ram_58__3)
          , .B1 (nx64920)) ;
    dffr reg_ram_59__3 (.Q (ram_59__3), .QB (\$dummy [874]), .D (nx42790), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42791 (.Y (nx42790), .A0 (ram_59__3), .A1 (nx65784), .S0 (nx63950
             )) ;
    dffr reg_ram_58__3 (.Q (ram_58__3), .QB (\$dummy [875]), .D (nx42800), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42801 (.Y (nx42800), .A0 (ram_58__3), .A1 (nx65784), .S0 (nx63954
             )) ;
    aoi22 ix58266 (.Y (nx58265), .A0 (ram_60__3), .A1 (nx64958), .B0 (ram_61__3)
          , .B1 (nx64996)) ;
    dffr reg_ram_60__3 (.Q (ram_60__3), .QB (\$dummy [876]), .D (nx42780), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42781 (.Y (nx42780), .A0 (ram_60__3), .A1 (nx65784), .S0 (nx63946
             )) ;
    dffr reg_ram_61__3 (.Q (ram_61__3), .QB (\$dummy [877]), .D (nx42770), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42771 (.Y (nx42770), .A0 (ram_61__3), .A1 (nx65784), .S0 (nx63942
             )) ;
    aoi22 ix58274 (.Y (nx58273), .A0 (ram_63__3), .A1 (nx65034), .B0 (ram_62__3)
          , .B1 (nx65072)) ;
    dffr reg_ram_63__3 (.Q (ram_63__3), .QB (\$dummy [878]), .D (nx42750), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42751 (.Y (nx42750), .A0 (ram_63__3), .A1 (nx65784), .S0 (nx63934
             )) ;
    dffr reg_ram_62__3 (.Q (ram_62__3), .QB (\$dummy [879]), .D (nx42760), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42761 (.Y (nx42760), .A0 (ram_62__3), .A1 (nx65784), .S0 (nx63938
             )) ;
    oai21 ix58282 (.Y (nx58281), .A0 (nx11506), .A1 (nx11428), .B0 (nx65124)) ;
    nand04 ix11507 (.Y (nx11506), .A0 (nx58284), .A1 (nx58292), .A2 (nx58300), .A3 (
           nx58308)) ;
    aoi22 ix58285 (.Y (nx58284), .A0 (ram_32__3), .A1 (nx64504), .B0 (ram_33__3)
          , .B1 (nx64542)) ;
    dffr reg_ram_32__3 (.Q (ram_32__3), .QB (\$dummy [880]), .D (nx42740), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42741 (.Y (nx42740), .A0 (ram_32__3), .A1 (nx65786), .S0 (nx63924
             )) ;
    dffr reg_ram_33__3 (.Q (ram_33__3), .QB (\$dummy [881]), .D (nx42730), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42731 (.Y (nx42730), .A0 (ram_33__3), .A1 (nx65786), .S0 (nx63920
             )) ;
    aoi22 ix58293 (.Y (nx58292), .A0 (ram_35__3), .A1 (nx64580), .B0 (ram_34__3)
          , .B1 (nx64618)) ;
    dffr reg_ram_35__3 (.Q (ram_35__3), .QB (\$dummy [882]), .D (nx42710), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42711 (.Y (nx42710), .A0 (ram_35__3), .A1 (nx65786), .S0 (nx63912
             )) ;
    dffr reg_ram_34__3 (.Q (ram_34__3), .QB (\$dummy [883]), .D (nx42720), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42721 (.Y (nx42720), .A0 (ram_34__3), .A1 (nx65786), .S0 (nx63916
             )) ;
    aoi22 ix58301 (.Y (nx58300), .A0 (ram_36__3), .A1 (nx64656), .B0 (ram_37__3)
          , .B1 (nx64694)) ;
    dffr reg_ram_36__3 (.Q (ram_36__3), .QB (\$dummy [884]), .D (nx42700), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42701 (.Y (nx42700), .A0 (ram_36__3), .A1 (nx65786), .S0 (nx63908
             )) ;
    dffr reg_ram_37__3 (.Q (ram_37__3), .QB (\$dummy [885]), .D (nx42690), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42691 (.Y (nx42690), .A0 (ram_37__3), .A1 (nx65786), .S0 (nx63904
             )) ;
    aoi22 ix58309 (.Y (nx58308), .A0 (ram_39__3), .A1 (nx64732), .B0 (ram_38__3)
          , .B1 (nx64770)) ;
    dffr reg_ram_39__3 (.Q (ram_39__3), .QB (\$dummy [886]), .D (nx42670), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42671 (.Y (nx42670), .A0 (ram_39__3), .A1 (nx65786), .S0 (nx63896
             )) ;
    dffr reg_ram_38__3 (.Q (ram_38__3), .QB (\$dummy [887]), .D (nx42680), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42681 (.Y (nx42680), .A0 (ram_38__3), .A1 (nx65788), .S0 (nx63900
             )) ;
    nand04 ix11429 (.Y (nx11428), .A0 (nx58317), .A1 (nx58325), .A2 (nx58333), .A3 (
           nx58341)) ;
    aoi22 ix58318 (.Y (nx58317), .A0 (ram_40__3), .A1 (nx64808), .B0 (ram_41__3)
          , .B1 (nx64846)) ;
    dffr reg_ram_40__3 (.Q (ram_40__3), .QB (\$dummy [888]), .D (nx42660), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42661 (.Y (nx42660), .A0 (ram_40__3), .A1 (nx65788), .S0 (nx63892
             )) ;
    dffr reg_ram_41__3 (.Q (ram_41__3), .QB (\$dummy [889]), .D (nx42650), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42651 (.Y (nx42650), .A0 (ram_41__3), .A1 (nx65788), .S0 (nx63888
             )) ;
    aoi22 ix58326 (.Y (nx58325), .A0 (ram_43__3), .A1 (nx64884), .B0 (ram_42__3)
          , .B1 (nx64922)) ;
    dffr reg_ram_43__3 (.Q (ram_43__3), .QB (\$dummy [890]), .D (nx42630), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42631 (.Y (nx42630), .A0 (ram_43__3), .A1 (nx65788), .S0 (nx63880
             )) ;
    dffr reg_ram_42__3 (.Q (ram_42__3), .QB (\$dummy [891]), .D (nx42640), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42641 (.Y (nx42640), .A0 (ram_42__3), .A1 (nx65788), .S0 (nx63884
             )) ;
    aoi22 ix58334 (.Y (nx58333), .A0 (ram_44__3), .A1 (nx64960), .B0 (ram_45__3)
          , .B1 (nx64998)) ;
    dffr reg_ram_44__3 (.Q (ram_44__3), .QB (\$dummy [892]), .D (nx42620), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42621 (.Y (nx42620), .A0 (ram_44__3), .A1 (nx65788), .S0 (nx63876
             )) ;
    dffr reg_ram_45__3 (.Q (ram_45__3), .QB (\$dummy [893]), .D (nx42610), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42611 (.Y (nx42610), .A0 (ram_45__3), .A1 (nx65788), .S0 (nx63872
             )) ;
    aoi22 ix58342 (.Y (nx58341), .A0 (ram_47__3), .A1 (nx65036), .B0 (ram_46__3)
          , .B1 (nx65074)) ;
    dffr reg_ram_47__3 (.Q (ram_47__3), .QB (\$dummy [894]), .D (nx42590), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42591 (.Y (nx42590), .A0 (ram_47__3), .A1 (nx65790), .S0 (nx63864
             )) ;
    dffr reg_ram_46__3 (.Q (ram_46__3), .QB (\$dummy [895]), .D (nx42600), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42601 (.Y (nx42600), .A0 (ram_46__3), .A1 (nx65790), .S0 (nx63868
             )) ;
    nand04 ix11349 (.Y (nx11348), .A0 (nx58350), .A1 (nx58418), .A2 (nx58486), .A3 (
           nx58554)) ;
    oai21 ix58351 (.Y (nx58350), .A0 (nx11338), .A1 (nx11260), .B0 (nx65128)) ;
    nand04 ix11339 (.Y (nx11338), .A0 (nx58353), .A1 (nx58361), .A2 (nx58369), .A3 (
           nx58377)) ;
    aoi22 ix58354 (.Y (nx58353), .A0 (ram_16__3), .A1 (nx64504), .B0 (ram_17__3)
          , .B1 (nx64542)) ;
    dffr reg_ram_16__3 (.Q (ram_16__3), .QB (\$dummy [896]), .D (nx42580), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42581 (.Y (nx42580), .A0 (ram_16__3), .A1 (nx65790), .S0 (nx63854
             )) ;
    dffr reg_ram_17__3 (.Q (ram_17__3), .QB (\$dummy [897]), .D (nx42570), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42571 (.Y (nx42570), .A0 (ram_17__3), .A1 (nx65790), .S0 (nx63850
             )) ;
    aoi22 ix58362 (.Y (nx58361), .A0 (ram_19__3), .A1 (nx64580), .B0 (ram_18__3)
          , .B1 (nx64618)) ;
    dffr reg_ram_19__3 (.Q (ram_19__3), .QB (\$dummy [898]), .D (nx42550), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42551 (.Y (nx42550), .A0 (ram_19__3), .A1 (nx65790), .S0 (nx63842
             )) ;
    dffr reg_ram_18__3 (.Q (ram_18__3), .QB (\$dummy [899]), .D (nx42560), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42561 (.Y (nx42560), .A0 (ram_18__3), .A1 (nx65790), .S0 (nx63846
             )) ;
    aoi22 ix58370 (.Y (nx58369), .A0 (ram_20__3), .A1 (nx64656), .B0 (ram_21__3)
          , .B1 (nx64694)) ;
    dffr reg_ram_20__3 (.Q (ram_20__3), .QB (\$dummy [900]), .D (nx42540), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42541 (.Y (nx42540), .A0 (ram_20__3), .A1 (nx65790), .S0 (nx63838
             )) ;
    dffr reg_ram_21__3 (.Q (ram_21__3), .QB (\$dummy [901]), .D (nx42530), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42531 (.Y (nx42530), .A0 (ram_21__3), .A1 (nx65792), .S0 (nx63834
             )) ;
    aoi22 ix58378 (.Y (nx58377), .A0 (ram_23__3), .A1 (nx64732), .B0 (ram_22__3)
          , .B1 (nx64770)) ;
    dffr reg_ram_23__3 (.Q (ram_23__3), .QB (\$dummy [902]), .D (nx42510), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42511 (.Y (nx42510), .A0 (ram_23__3), .A1 (nx65792), .S0 (nx63826
             )) ;
    dffr reg_ram_22__3 (.Q (ram_22__3), .QB (\$dummy [903]), .D (nx42520), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42521 (.Y (nx42520), .A0 (ram_22__3), .A1 (nx65792), .S0 (nx63830
             )) ;
    nand04 ix11261 (.Y (nx11260), .A0 (nx58386), .A1 (nx58394), .A2 (nx58402), .A3 (
           nx58410)) ;
    aoi22 ix58387 (.Y (nx58386), .A0 (ram_24__3), .A1 (nx64808), .B0 (ram_25__3)
          , .B1 (nx64846)) ;
    dffr reg_ram_24__3 (.Q (ram_24__3), .QB (\$dummy [904]), .D (nx42500), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42501 (.Y (nx42500), .A0 (ram_24__3), .A1 (nx65792), .S0 (nx63822
             )) ;
    dffr reg_ram_25__3 (.Q (ram_25__3), .QB (\$dummy [905]), .D (nx42490), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42491 (.Y (nx42490), .A0 (ram_25__3), .A1 (nx65792), .S0 (nx63818
             )) ;
    aoi22 ix58395 (.Y (nx58394), .A0 (ram_27__3), .A1 (nx64884), .B0 (ram_26__3)
          , .B1 (nx64922)) ;
    dffr reg_ram_27__3 (.Q (ram_27__3), .QB (\$dummy [906]), .D (nx42470), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42471 (.Y (nx42470), .A0 (ram_27__3), .A1 (nx65792), .S0 (nx63810
             )) ;
    dffr reg_ram_26__3 (.Q (ram_26__3), .QB (\$dummy [907]), .D (nx42480), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42481 (.Y (nx42480), .A0 (ram_26__3), .A1 (nx65792), .S0 (nx63814
             )) ;
    aoi22 ix58403 (.Y (nx58402), .A0 (ram_28__3), .A1 (nx64960), .B0 (ram_29__3)
          , .B1 (nx64998)) ;
    dffr reg_ram_28__3 (.Q (ram_28__3), .QB (\$dummy [908]), .D (nx42460), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42461 (.Y (nx42460), .A0 (ram_28__3), .A1 (nx65794), .S0 (nx63806
             )) ;
    dffr reg_ram_29__3 (.Q (ram_29__3), .QB (\$dummy [909]), .D (nx42450), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42451 (.Y (nx42450), .A0 (ram_29__3), .A1 (nx65794), .S0 (nx63802
             )) ;
    aoi22 ix58411 (.Y (nx58410), .A0 (ram_31__3), .A1 (nx65036), .B0 (ram_30__3)
          , .B1 (nx65074)) ;
    dffr reg_ram_31__3 (.Q (ram_31__3), .QB (\$dummy [910]), .D (nx42430), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42431 (.Y (nx42430), .A0 (ram_31__3), .A1 (nx65794), .S0 (nx63794
             )) ;
    dffr reg_ram_30__3 (.Q (ram_30__3), .QB (\$dummy [911]), .D (nx42440), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42441 (.Y (nx42440), .A0 (ram_30__3), .A1 (nx65794), .S0 (nx63798
             )) ;
    oai21 ix58419 (.Y (nx58418), .A0 (nx11176), .A1 (nx11098), .B0 (nx65142)) ;
    nand04 ix11177 (.Y (nx11176), .A0 (nx58421), .A1 (nx58429), .A2 (nx58437), .A3 (
           nx58445)) ;
    aoi22 ix58422 (.Y (nx58421), .A0 (ram_0__3), .A1 (nx64504), .B0 (ram_1__3), 
          .B1 (nx64542)) ;
    dffr reg_ram_0__3 (.Q (ram_0__3), .QB (\$dummy [912]), .D (nx42420), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42421 (.Y (nx42420), .A0 (nx65794), .A1 (ram_0__3), .S0 (nx65132)
             ) ;
    dffr reg_ram_1__3 (.Q (ram_1__3), .QB (\$dummy [913]), .D (nx42410), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42411 (.Y (nx42410), .A0 (nx65794), .A1 (ram_1__3), .S0 (nx65146)
             ) ;
    aoi22 ix58430 (.Y (nx58429), .A0 (ram_3__3), .A1 (nx64580), .B0 (ram_2__3), 
          .B1 (nx64618)) ;
    dffr reg_ram_3__3 (.Q (ram_3__3), .QB (\$dummy [914]), .D (nx42390), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42391 (.Y (nx42390), .A0 (nx65794), .A1 (ram_3__3), .S0 (nx65150)
             ) ;
    dffr reg_ram_2__3 (.Q (ram_2__3), .QB (\$dummy [915]), .D (nx42400), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42401 (.Y (nx42400), .A0 (nx65796), .A1 (ram_2__3), .S0 (nx65154)
             ) ;
    aoi22 ix58438 (.Y (nx58437), .A0 (ram_4__3), .A1 (nx64656), .B0 (ram_5__3), 
          .B1 (nx64694)) ;
    dffr reg_ram_4__3 (.Q (ram_4__3), .QB (\$dummy [916]), .D (nx42380), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42381 (.Y (nx42380), .A0 (nx65796), .A1 (ram_4__3), .S0 (nx65158)
             ) ;
    dffr reg_ram_5__3 (.Q (ram_5__3), .QB (\$dummy [917]), .D (nx42370), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42371 (.Y (nx42370), .A0 (nx65796), .A1 (ram_5__3), .S0 (nx65162)
             ) ;
    aoi22 ix58446 (.Y (nx58445), .A0 (ram_7__3), .A1 (nx64732), .B0 (ram_6__3), 
          .B1 (nx64770)) ;
    dffr reg_ram_7__3 (.Q (ram_7__3), .QB (\$dummy [918]), .D (nx42350), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42351 (.Y (nx42350), .A0 (nx65796), .A1 (ram_7__3), .S0 (nx65166)
             ) ;
    dffr reg_ram_6__3 (.Q (ram_6__3), .QB (\$dummy [919]), .D (nx42360), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42361 (.Y (nx42360), .A0 (nx65796), .A1 (ram_6__3), .S0 (nx65170)
             ) ;
    nand04 ix11099 (.Y (nx11098), .A0 (nx58454), .A1 (nx58462), .A2 (nx58470), .A3 (
           nx58478)) ;
    aoi22 ix58455 (.Y (nx58454), .A0 (ram_8__3), .A1 (nx64808), .B0 (ram_9__3), 
          .B1 (nx64846)) ;
    dffr reg_ram_8__3 (.Q (ram_8__3), .QB (\$dummy [920]), .D (nx42340), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42341 (.Y (nx42340), .A0 (nx65796), .A1 (ram_8__3), .S0 (nx65174)
             ) ;
    dffr reg_ram_9__3 (.Q (ram_9__3), .QB (\$dummy [921]), .D (nx42330), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42331 (.Y (nx42330), .A0 (nx65796), .A1 (ram_9__3), .S0 (nx65178)
             ) ;
    aoi22 ix58463 (.Y (nx58462), .A0 (ram_11__3), .A1 (nx64884), .B0 (ram_10__3)
          , .B1 (nx64922)) ;
    dffr reg_ram_11__3 (.Q (ram_11__3), .QB (\$dummy [922]), .D (nx42310), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42311 (.Y (nx42310), .A0 (nx65798), .A1 (ram_11__3), .S0 (nx65182
             )) ;
    dffr reg_ram_10__3 (.Q (ram_10__3), .QB (\$dummy [923]), .D (nx42320), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42321 (.Y (nx42320), .A0 (nx65798), .A1 (ram_10__3), .S0 (nx65186
             )) ;
    aoi22 ix58471 (.Y (nx58470), .A0 (ram_12__3), .A1 (nx64960), .B0 (ram_13__3)
          , .B1 (nx64998)) ;
    dffr reg_ram_12__3 (.Q (ram_12__3), .QB (\$dummy [924]), .D (nx42300), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42301 (.Y (nx42300), .A0 (nx65798), .A1 (ram_12__3), .S0 (nx65190
             )) ;
    dffr reg_ram_13__3 (.Q (ram_13__3), .QB (\$dummy [925]), .D (nx42290), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42291 (.Y (nx42290), .A0 (nx65798), .A1 (ram_13__3), .S0 (nx65194
             )) ;
    aoi22 ix58479 (.Y (nx58478), .A0 (ram_15__3), .A1 (nx65036), .B0 (ram_14__3)
          , .B1 (nx65074)) ;
    dffr reg_ram_15__3 (.Q (ram_15__3), .QB (\$dummy [926]), .D (nx42270), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42271 (.Y (nx42270), .A0 (nx65798), .A1 (ram_15__3), .S0 (nx65198
             )) ;
    dffr reg_ram_14__3 (.Q (ram_14__3), .QB (\$dummy [927]), .D (nx42280), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42281 (.Y (nx42280), .A0 (nx65798), .A1 (ram_14__3), .S0 (nx65202
             )) ;
    oai21 ix58487 (.Y (nx58486), .A0 (nx11012), .A1 (nx10934), .B0 (nx65206)) ;
    nand04 ix11013 (.Y (nx11012), .A0 (nx58489), .A1 (nx58497), .A2 (nx58505), .A3 (
           nx58513)) ;
    aoi22 ix58490 (.Y (nx58489), .A0 (ram_96__3), .A1 (nx64504), .B0 (ram_97__3)
          , .B1 (nx64542)) ;
    dffr reg_ram_96__3 (.Q (ram_96__3), .QB (\$dummy [928]), .D (nx42260), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42261 (.Y (nx42260), .A0 (ram_96__3), .A1 (nx65798), .S0 (nx63784
             )) ;
    dffr reg_ram_97__3 (.Q (ram_97__3), .QB (\$dummy [929]), .D (nx42250), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42251 (.Y (nx42250), .A0 (ram_97__3), .A1 (nx65800), .S0 (nx63780
             )) ;
    aoi22 ix58498 (.Y (nx58497), .A0 (ram_99__3), .A1 (nx64580), .B0 (ram_98__3)
          , .B1 (nx64618)) ;
    dffr reg_ram_99__3 (.Q (ram_99__3), .QB (\$dummy [930]), .D (nx42230), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42231 (.Y (nx42230), .A0 (ram_99__3), .A1 (nx65800), .S0 (nx63772
             )) ;
    dffr reg_ram_98__3 (.Q (ram_98__3), .QB (\$dummy [931]), .D (nx42240), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42241 (.Y (nx42240), .A0 (ram_98__3), .A1 (nx65800), .S0 (nx63776
             )) ;
    aoi22 ix58506 (.Y (nx58505), .A0 (ram_100__3), .A1 (nx64656), .B0 (
          ram_101__3), .B1 (nx64694)) ;
    dffr reg_ram_100__3 (.Q (ram_100__3), .QB (\$dummy [932]), .D (nx42220), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42221 (.Y (nx42220), .A0 (ram_100__3), .A1 (nx65800), .S0 (
             nx63768)) ;
    dffr reg_ram_101__3 (.Q (ram_101__3), .QB (\$dummy [933]), .D (nx42210), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42211 (.Y (nx42210), .A0 (ram_101__3), .A1 (nx65800), .S0 (
             nx63764)) ;
    aoi22 ix58514 (.Y (nx58513), .A0 (ram_103__3), .A1 (nx64732), .B0 (
          ram_102__3), .B1 (nx64770)) ;
    dffr reg_ram_103__3 (.Q (ram_103__3), .QB (\$dummy [934]), .D (nx42190), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42191 (.Y (nx42190), .A0 (ram_103__3), .A1 (nx65800), .S0 (
             nx63756)) ;
    dffr reg_ram_102__3 (.Q (ram_102__3), .QB (\$dummy [935]), .D (nx42200), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42201 (.Y (nx42200), .A0 (ram_102__3), .A1 (nx65800), .S0 (
             nx63760)) ;
    nand04 ix10935 (.Y (nx10934), .A0 (nx58522), .A1 (nx58530), .A2 (nx58538), .A3 (
           nx58546)) ;
    aoi22 ix58523 (.Y (nx58522), .A0 (ram_104__3), .A1 (nx64808), .B0 (
          ram_105__3), .B1 (nx64846)) ;
    dffr reg_ram_104__3 (.Q (ram_104__3), .QB (\$dummy [936]), .D (nx42180), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42181 (.Y (nx42180), .A0 (ram_104__3), .A1 (nx65802), .S0 (
             nx63752)) ;
    dffr reg_ram_105__3 (.Q (ram_105__3), .QB (\$dummy [937]), .D (nx42170), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42171 (.Y (nx42170), .A0 (ram_105__3), .A1 (nx65802), .S0 (
             nx63748)) ;
    aoi22 ix58531 (.Y (nx58530), .A0 (ram_107__3), .A1 (nx64884), .B0 (
          ram_106__3), .B1 (nx64922)) ;
    dffr reg_ram_107__3 (.Q (ram_107__3), .QB (\$dummy [938]), .D (nx42150), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42151 (.Y (nx42150), .A0 (ram_107__3), .A1 (nx65802), .S0 (
             nx63740)) ;
    dffr reg_ram_106__3 (.Q (ram_106__3), .QB (\$dummy [939]), .D (nx42160), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42161 (.Y (nx42160), .A0 (ram_106__3), .A1 (nx65802), .S0 (
             nx63744)) ;
    aoi22 ix58539 (.Y (nx58538), .A0 (ram_108__3), .A1 (nx64960), .B0 (
          ram_109__3), .B1 (nx64998)) ;
    dffr reg_ram_108__3 (.Q (ram_108__3), .QB (\$dummy [940]), .D (nx42140), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42141 (.Y (nx42140), .A0 (ram_108__3), .A1 (nx65802), .S0 (
             nx63736)) ;
    dffr reg_ram_109__3 (.Q (ram_109__3), .QB (\$dummy [941]), .D (nx42130), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42131 (.Y (nx42130), .A0 (ram_109__3), .A1 (nx65802), .S0 (
             nx63732)) ;
    aoi22 ix58547 (.Y (nx58546), .A0 (ram_111__3), .A1 (nx65036), .B0 (
          ram_110__3), .B1 (nx65074)) ;
    dffr reg_ram_111__3 (.Q (ram_111__3), .QB (\$dummy [942]), .D (nx42110), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42111 (.Y (nx42110), .A0 (ram_111__3), .A1 (nx65802), .S0 (
             nx63724)) ;
    dffr reg_ram_110__3 (.Q (ram_110__3), .QB (\$dummy [943]), .D (nx42120), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42121 (.Y (nx42120), .A0 (ram_110__3), .A1 (nx65804), .S0 (
             nx63728)) ;
    oai21 ix58555 (.Y (nx58554), .A0 (nx10850), .A1 (nx10772), .B0 (nx65210)) ;
    nand04 ix10851 (.Y (nx10850), .A0 (nx58557), .A1 (nx58565), .A2 (nx58573), .A3 (
           nx58581)) ;
    aoi22 ix58558 (.Y (nx58557), .A0 (ram_112__3), .A1 (nx64504), .B0 (
          ram_113__3), .B1 (nx64542)) ;
    dffr reg_ram_112__3 (.Q (ram_112__3), .QB (\$dummy [944]), .D (nx42100), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42101 (.Y (nx42100), .A0 (ram_112__3), .A1 (nx65804), .S0 (
             nx63714)) ;
    dffr reg_ram_113__3 (.Q (ram_113__3), .QB (\$dummy [945]), .D (nx42090), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42091 (.Y (nx42090), .A0 (ram_113__3), .A1 (nx65804), .S0 (
             nx63710)) ;
    aoi22 ix58566 (.Y (nx58565), .A0 (ram_115__3), .A1 (nx64580), .B0 (
          ram_114__3), .B1 (nx64618)) ;
    dffr reg_ram_115__3 (.Q (ram_115__3), .QB (\$dummy [946]), .D (nx42070), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42071 (.Y (nx42070), .A0 (ram_115__3), .A1 (nx65804), .S0 (
             nx63702)) ;
    dffr reg_ram_114__3 (.Q (ram_114__3), .QB (\$dummy [947]), .D (nx42080), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42081 (.Y (nx42080), .A0 (ram_114__3), .A1 (nx65804), .S0 (
             nx63706)) ;
    aoi22 ix58574 (.Y (nx58573), .A0 (ram_116__3), .A1 (nx64656), .B0 (
          ram_117__3), .B1 (nx64694)) ;
    dffr reg_ram_116__3 (.Q (ram_116__3), .QB (\$dummy [948]), .D (nx42060), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42061 (.Y (nx42060), .A0 (ram_116__3), .A1 (nx65804), .S0 (
             nx63698)) ;
    dffr reg_ram_117__3 (.Q (ram_117__3), .QB (\$dummy [949]), .D (nx42050), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42051 (.Y (nx42050), .A0 (ram_117__3), .A1 (nx65804), .S0 (
             nx63694)) ;
    aoi22 ix58582 (.Y (nx58581), .A0 (ram_119__3), .A1 (nx64732), .B0 (
          ram_118__3), .B1 (nx64770)) ;
    dffr reg_ram_119__3 (.Q (ram_119__3), .QB (\$dummy [950]), .D (nx42030), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42031 (.Y (nx42030), .A0 (ram_119__3), .A1 (nx65806), .S0 (
             nx63686)) ;
    dffr reg_ram_118__3 (.Q (ram_118__3), .QB (\$dummy [951]), .D (nx42040), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42041 (.Y (nx42040), .A0 (ram_118__3), .A1 (nx65806), .S0 (
             nx63690)) ;
    nand04 ix10773 (.Y (nx10772), .A0 (nx58590), .A1 (nx58598), .A2 (nx58606), .A3 (
           nx58614)) ;
    aoi22 ix58591 (.Y (nx58590), .A0 (ram_120__3), .A1 (nx64808), .B0 (
          ram_121__3), .B1 (nx64846)) ;
    dffr reg_ram_120__3 (.Q (ram_120__3), .QB (\$dummy [952]), .D (nx42020), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42021 (.Y (nx42020), .A0 (ram_120__3), .A1 (nx65806), .S0 (
             nx63682)) ;
    dffr reg_ram_121__3 (.Q (ram_121__3), .QB (\$dummy [953]), .D (nx42010), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42011 (.Y (nx42010), .A0 (ram_121__3), .A1 (nx65806), .S0 (
             nx63678)) ;
    aoi22 ix58599 (.Y (nx58598), .A0 (ram_123__3), .A1 (nx64884), .B0 (
          ram_122__3), .B1 (nx64922)) ;
    dffr reg_ram_123__3 (.Q (ram_123__3), .QB (\$dummy [954]), .D (nx41990), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41991 (.Y (nx41990), .A0 (ram_123__3), .A1 (nx65806), .S0 (
             nx63670)) ;
    dffr reg_ram_122__3 (.Q (ram_122__3), .QB (\$dummy [955]), .D (nx42000), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix42001 (.Y (nx42000), .A0 (ram_122__3), .A1 (nx65806), .S0 (
             nx63674)) ;
    aoi22 ix58607 (.Y (nx58606), .A0 (ram_124__3), .A1 (nx64960), .B0 (
          ram_125__3), .B1 (nx64998)) ;
    dffr reg_ram_124__3 (.Q (ram_124__3), .QB (\$dummy [956]), .D (nx41980), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41981 (.Y (nx41980), .A0 (ram_124__3), .A1 (nx65806), .S0 (
             nx63666)) ;
    dffr reg_ram_125__3 (.Q (ram_125__3), .QB (\$dummy [957]), .D (nx41970), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41971 (.Y (nx41970), .A0 (ram_125__3), .A1 (nx65808), .S0 (
             nx63662)) ;
    aoi22 ix58615 (.Y (nx58614), .A0 (ram_127__3), .A1 (nx65036), .B0 (
          ram_126__3), .B1 (nx65074)) ;
    dffr reg_ram_127__3 (.Q (ram_127__3), .QB (\$dummy [958]), .D (nx41950), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41951 (.Y (nx41950), .A0 (ram_127__3), .A1 (nx65808), .S0 (
             nx63654)) ;
    dffr reg_ram_126__3 (.Q (ram_126__3), .QB (\$dummy [959]), .D (nx41960), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41961 (.Y (nx41960), .A0 (ram_126__3), .A1 (nx65808), .S0 (
             nx63658)) ;
    nand04 ix10695 (.Y (nx10694), .A0 (nx58623), .A1 (nx58691), .A2 (nx58759), .A3 (
           nx58827)) ;
    oai21 ix58624 (.Y (nx58623), .A0 (nx10684), .A1 (nx10606), .B0 (nx65214)) ;
    nand04 ix10685 (.Y (nx10684), .A0 (nx58626), .A1 (nx58634), .A2 (nx58642), .A3 (
           nx58650)) ;
    aoi22 ix58627 (.Y (nx58626), .A0 (ram_128__3), .A1 (nx64504), .B0 (
          ram_129__3), .B1 (nx64542)) ;
    dffr reg_ram_128__3 (.Q (ram_128__3), .QB (\$dummy [960]), .D (nx41940), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41941 (.Y (nx41940), .A0 (ram_128__3), .A1 (nx65808), .S0 (
             nx63644)) ;
    dffr reg_ram_129__3 (.Q (ram_129__3), .QB (\$dummy [961]), .D (nx41930), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41931 (.Y (nx41930), .A0 (ram_129__3), .A1 (nx65808), .S0 (
             nx63640)) ;
    aoi22 ix58635 (.Y (nx58634), .A0 (ram_131__3), .A1 (nx64580), .B0 (
          ram_130__3), .B1 (nx64618)) ;
    dffr reg_ram_131__3 (.Q (ram_131__3), .QB (\$dummy [962]), .D (nx41910), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41911 (.Y (nx41910), .A0 (ram_131__3), .A1 (nx65808), .S0 (
             nx63632)) ;
    dffr reg_ram_130__3 (.Q (ram_130__3), .QB (\$dummy [963]), .D (nx41920), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41921 (.Y (nx41920), .A0 (ram_130__3), .A1 (nx65808), .S0 (
             nx63636)) ;
    aoi22 ix58643 (.Y (nx58642), .A0 (ram_132__3), .A1 (nx64656), .B0 (
          ram_133__3), .B1 (nx64694)) ;
    dffr reg_ram_132__3 (.Q (ram_132__3), .QB (\$dummy [964]), .D (nx41900), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41901 (.Y (nx41900), .A0 (ram_132__3), .A1 (nx65810), .S0 (
             nx63628)) ;
    dffr reg_ram_133__3 (.Q (ram_133__3), .QB (\$dummy [965]), .D (nx41890), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41891 (.Y (nx41890), .A0 (ram_133__3), .A1 (nx65810), .S0 (
             nx63624)) ;
    aoi22 ix58651 (.Y (nx58650), .A0 (ram_135__3), .A1 (nx64732), .B0 (
          ram_134__3), .B1 (nx64770)) ;
    dffr reg_ram_135__3 (.Q (ram_135__3), .QB (\$dummy [966]), .D (nx41870), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41871 (.Y (nx41870), .A0 (ram_135__3), .A1 (nx65810), .S0 (
             nx63616)) ;
    dffr reg_ram_134__3 (.Q (ram_134__3), .QB (\$dummy [967]), .D (nx41880), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41881 (.Y (nx41880), .A0 (ram_134__3), .A1 (nx65810), .S0 (
             nx63620)) ;
    nand04 ix10607 (.Y (nx10606), .A0 (nx58659), .A1 (nx58667), .A2 (nx58675), .A3 (
           nx58683)) ;
    aoi22 ix58660 (.Y (nx58659), .A0 (ram_136__3), .A1 (nx64808), .B0 (
          ram_137__3), .B1 (nx64846)) ;
    dffr reg_ram_136__3 (.Q (ram_136__3), .QB (\$dummy [968]), .D (nx41860), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41861 (.Y (nx41860), .A0 (ram_136__3), .A1 (nx65810), .S0 (
             nx63612)) ;
    dffr reg_ram_137__3 (.Q (ram_137__3), .QB (\$dummy [969]), .D (nx41850), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41851 (.Y (nx41850), .A0 (ram_137__3), .A1 (nx65810), .S0 (
             nx63608)) ;
    aoi22 ix58668 (.Y (nx58667), .A0 (ram_139__3), .A1 (nx64884), .B0 (
          ram_138__3), .B1 (nx64922)) ;
    dffr reg_ram_139__3 (.Q (ram_139__3), .QB (\$dummy [970]), .D (nx41830), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41831 (.Y (nx41830), .A0 (ram_139__3), .A1 (nx65810), .S0 (
             nx63600)) ;
    dffr reg_ram_138__3 (.Q (ram_138__3), .QB (\$dummy [971]), .D (nx41840), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41841 (.Y (nx41840), .A0 (ram_138__3), .A1 (nx65812), .S0 (
             nx63604)) ;
    aoi22 ix58676 (.Y (nx58675), .A0 (ram_140__3), .A1 (nx64960), .B0 (
          ram_141__3), .B1 (nx64998)) ;
    dffr reg_ram_140__3 (.Q (ram_140__3), .QB (\$dummy [972]), .D (nx41820), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41821 (.Y (nx41820), .A0 (ram_140__3), .A1 (nx65812), .S0 (
             nx63596)) ;
    dffr reg_ram_141__3 (.Q (ram_141__3), .QB (\$dummy [973]), .D (nx41810), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41811 (.Y (nx41810), .A0 (ram_141__3), .A1 (nx65812), .S0 (
             nx63592)) ;
    aoi22 ix58684 (.Y (nx58683), .A0 (ram_143__3), .A1 (nx65036), .B0 (
          ram_142__3), .B1 (nx65074)) ;
    dffr reg_ram_143__3 (.Q (ram_143__3), .QB (\$dummy [974]), .D (nx41790), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41791 (.Y (nx41790), .A0 (ram_143__3), .A1 (nx65812), .S0 (
             nx63584)) ;
    dffr reg_ram_142__3 (.Q (ram_142__3), .QB (\$dummy [975]), .D (nx41800), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41801 (.Y (nx41800), .A0 (ram_142__3), .A1 (nx65812), .S0 (
             nx63588)) ;
    oai21 ix58692 (.Y (nx58691), .A0 (nx10522), .A1 (nx10444), .B0 (nx65218)) ;
    nand04 ix10523 (.Y (nx10522), .A0 (nx58694), .A1 (nx58702), .A2 (nx58710), .A3 (
           nx58718)) ;
    aoi22 ix58695 (.Y (nx58694), .A0 (ram_144__3), .A1 (nx64504), .B0 (
          ram_145__3), .B1 (nx64542)) ;
    dffr reg_ram_144__3 (.Q (ram_144__3), .QB (\$dummy [976]), .D (nx41780), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41781 (.Y (nx41780), .A0 (ram_144__3), .A1 (nx65812), .S0 (
             nx63574)) ;
    dffr reg_ram_145__3 (.Q (ram_145__3), .QB (\$dummy [977]), .D (nx41770), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41771 (.Y (nx41770), .A0 (ram_145__3), .A1 (nx65812), .S0 (
             nx63570)) ;
    aoi22 ix58703 (.Y (nx58702), .A0 (ram_147__3), .A1 (nx64580), .B0 (
          ram_146__3), .B1 (nx64618)) ;
    dffr reg_ram_147__3 (.Q (ram_147__3), .QB (\$dummy [978]), .D (nx41750), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41751 (.Y (nx41750), .A0 (ram_147__3), .A1 (nx65814), .S0 (
             nx63562)) ;
    dffr reg_ram_146__3 (.Q (ram_146__3), .QB (\$dummy [979]), .D (nx41760), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41761 (.Y (nx41760), .A0 (ram_146__3), .A1 (nx65814), .S0 (
             nx63566)) ;
    aoi22 ix58711 (.Y (nx58710), .A0 (ram_148__3), .A1 (nx64656), .B0 (
          ram_149__3), .B1 (nx64694)) ;
    dffr reg_ram_148__3 (.Q (ram_148__3), .QB (\$dummy [980]), .D (nx41740), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41741 (.Y (nx41740), .A0 (ram_148__3), .A1 (nx65814), .S0 (
             nx63558)) ;
    dffr reg_ram_149__3 (.Q (ram_149__3), .QB (\$dummy [981]), .D (nx41730), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41731 (.Y (nx41730), .A0 (ram_149__3), .A1 (nx65814), .S0 (
             nx63554)) ;
    aoi22 ix58719 (.Y (nx58718), .A0 (ram_151__3), .A1 (nx64732), .B0 (
          ram_150__3), .B1 (nx64770)) ;
    dffr reg_ram_151__3 (.Q (ram_151__3), .QB (\$dummy [982]), .D (nx41710), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41711 (.Y (nx41710), .A0 (ram_151__3), .A1 (nx65814), .S0 (
             nx63546)) ;
    dffr reg_ram_150__3 (.Q (ram_150__3), .QB (\$dummy [983]), .D (nx41720), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41721 (.Y (nx41720), .A0 (ram_150__3), .A1 (nx65814), .S0 (
             nx63550)) ;
    nand04 ix10445 (.Y (nx10444), .A0 (nx58727), .A1 (nx58735), .A2 (nx58743), .A3 (
           nx58751)) ;
    aoi22 ix58728 (.Y (nx58727), .A0 (ram_152__3), .A1 (nx64808), .B0 (
          ram_153__3), .B1 (nx64846)) ;
    dffr reg_ram_152__3 (.Q (ram_152__3), .QB (\$dummy [984]), .D (nx41700), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41701 (.Y (nx41700), .A0 (ram_152__3), .A1 (nx65814), .S0 (
             nx63542)) ;
    dffr reg_ram_153__3 (.Q (ram_153__3), .QB (\$dummy [985]), .D (nx41690), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41691 (.Y (nx41690), .A0 (ram_153__3), .A1 (nx65816), .S0 (
             nx63538)) ;
    aoi22 ix58736 (.Y (nx58735), .A0 (ram_155__3), .A1 (nx64884), .B0 (
          ram_154__3), .B1 (nx64922)) ;
    dffr reg_ram_155__3 (.Q (ram_155__3), .QB (\$dummy [986]), .D (nx41670), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41671 (.Y (nx41670), .A0 (ram_155__3), .A1 (nx65816), .S0 (
             nx63530)) ;
    dffr reg_ram_154__3 (.Q (ram_154__3), .QB (\$dummy [987]), .D (nx41680), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41681 (.Y (nx41680), .A0 (ram_154__3), .A1 (nx65816), .S0 (
             nx63534)) ;
    aoi22 ix58744 (.Y (nx58743), .A0 (ram_156__3), .A1 (nx64960), .B0 (
          ram_157__3), .B1 (nx64998)) ;
    dffr reg_ram_156__3 (.Q (ram_156__3), .QB (\$dummy [988]), .D (nx41660), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41661 (.Y (nx41660), .A0 (ram_156__3), .A1 (nx65816), .S0 (
             nx63526)) ;
    dffr reg_ram_157__3 (.Q (ram_157__3), .QB (\$dummy [989]), .D (nx41650), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41651 (.Y (nx41650), .A0 (ram_157__3), .A1 (nx65816), .S0 (
             nx63522)) ;
    aoi22 ix58752 (.Y (nx58751), .A0 (ram_159__3), .A1 (nx65036), .B0 (
          ram_158__3), .B1 (nx65074)) ;
    dffr reg_ram_159__3 (.Q (ram_159__3), .QB (\$dummy [990]), .D (nx41630), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41631 (.Y (nx41630), .A0 (ram_159__3), .A1 (nx65816), .S0 (
             nx63514)) ;
    dffr reg_ram_158__3 (.Q (ram_158__3), .QB (\$dummy [991]), .D (nx41640), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41641 (.Y (nx41640), .A0 (ram_158__3), .A1 (nx65816), .S0 (
             nx63518)) ;
    oai21 ix58760 (.Y (nx58759), .A0 (nx10358), .A1 (nx10280), .B0 (nx65222)) ;
    nand04 ix10359 (.Y (nx10358), .A0 (nx58762), .A1 (nx58770), .A2 (nx58778), .A3 (
           nx58786)) ;
    aoi22 ix58763 (.Y (nx58762), .A0 (ram_160__3), .A1 (nx64506), .B0 (
          ram_161__3), .B1 (nx64544)) ;
    dffr reg_ram_160__3 (.Q (ram_160__3), .QB (\$dummy [992]), .D (nx41620), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41621 (.Y (nx41620), .A0 (ram_160__3), .A1 (nx65818), .S0 (
             nx63504)) ;
    dffr reg_ram_161__3 (.Q (ram_161__3), .QB (\$dummy [993]), .D (nx41610), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41611 (.Y (nx41610), .A0 (ram_161__3), .A1 (nx65818), .S0 (
             nx63500)) ;
    aoi22 ix58771 (.Y (nx58770), .A0 (ram_163__3), .A1 (nx64582), .B0 (
          ram_162__3), .B1 (nx64620)) ;
    dffr reg_ram_163__3 (.Q (ram_163__3), .QB (\$dummy [994]), .D (nx41590), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41591 (.Y (nx41590), .A0 (ram_163__3), .A1 (nx65818), .S0 (
             nx63492)) ;
    dffr reg_ram_162__3 (.Q (ram_162__3), .QB (\$dummy [995]), .D (nx41600), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41601 (.Y (nx41600), .A0 (ram_162__3), .A1 (nx65818), .S0 (
             nx63496)) ;
    aoi22 ix58779 (.Y (nx58778), .A0 (ram_164__3), .A1 (nx64658), .B0 (
          ram_165__3), .B1 (nx64696)) ;
    dffr reg_ram_164__3 (.Q (ram_164__3), .QB (\$dummy [996]), .D (nx41580), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41581 (.Y (nx41580), .A0 (ram_164__3), .A1 (nx65818), .S0 (
             nx63488)) ;
    dffr reg_ram_165__3 (.Q (ram_165__3), .QB (\$dummy [997]), .D (nx41570), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41571 (.Y (nx41570), .A0 (ram_165__3), .A1 (nx65818), .S0 (
             nx63484)) ;
    aoi22 ix58787 (.Y (nx58786), .A0 (ram_167__3), .A1 (nx64734), .B0 (
          ram_166__3), .B1 (nx64772)) ;
    dffr reg_ram_167__3 (.Q (ram_167__3), .QB (\$dummy [998]), .D (nx41550), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41551 (.Y (nx41550), .A0 (ram_167__3), .A1 (nx65818), .S0 (
             nx63476)) ;
    dffr reg_ram_166__3 (.Q (ram_166__3), .QB (\$dummy [999]), .D (nx41560), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41561 (.Y (nx41560), .A0 (ram_166__3), .A1 (nx65820), .S0 (
             nx63480)) ;
    nand04 ix10281 (.Y (nx10280), .A0 (nx58795), .A1 (nx58803), .A2 (nx58811), .A3 (
           nx58819)) ;
    aoi22 ix58796 (.Y (nx58795), .A0 (ram_168__3), .A1 (nx64810), .B0 (
          ram_169__3), .B1 (nx64848)) ;
    dffr reg_ram_168__3 (.Q (ram_168__3), .QB (\$dummy [1000]), .D (nx41540), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41541 (.Y (nx41540), .A0 (ram_168__3), .A1 (nx65820), .S0 (
             nx63472)) ;
    dffr reg_ram_169__3 (.Q (ram_169__3), .QB (\$dummy [1001]), .D (nx41530), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41531 (.Y (nx41530), .A0 (ram_169__3), .A1 (nx65820), .S0 (
             nx63468)) ;
    aoi22 ix58804 (.Y (nx58803), .A0 (ram_171__3), .A1 (nx64886), .B0 (
          ram_170__3), .B1 (nx64924)) ;
    dffr reg_ram_171__3 (.Q (ram_171__3), .QB (\$dummy [1002]), .D (nx41510), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41511 (.Y (nx41510), .A0 (ram_171__3), .A1 (nx65820), .S0 (
             nx63460)) ;
    dffr reg_ram_170__3 (.Q (ram_170__3), .QB (\$dummy [1003]), .D (nx41520), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41521 (.Y (nx41520), .A0 (ram_170__3), .A1 (nx65820), .S0 (
             nx63464)) ;
    aoi22 ix58812 (.Y (nx58811), .A0 (ram_172__3), .A1 (nx64962), .B0 (
          ram_173__3), .B1 (nx65000)) ;
    dffr reg_ram_172__3 (.Q (ram_172__3), .QB (\$dummy [1004]), .D (nx41500), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41501 (.Y (nx41500), .A0 (ram_172__3), .A1 (nx65820), .S0 (
             nx63456)) ;
    dffr reg_ram_173__3 (.Q (ram_173__3), .QB (\$dummy [1005]), .D (nx41490), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41491 (.Y (nx41490), .A0 (ram_173__3), .A1 (nx65820), .S0 (
             nx63452)) ;
    aoi22 ix58820 (.Y (nx58819), .A0 (ram_175__3), .A1 (nx65038), .B0 (
          ram_174__3), .B1 (nx65076)) ;
    dffr reg_ram_175__3 (.Q (ram_175__3), .QB (\$dummy [1006]), .D (nx41470), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41471 (.Y (nx41470), .A0 (ram_175__3), .A1 (nx65822), .S0 (
             nx63444)) ;
    dffr reg_ram_174__3 (.Q (ram_174__3), .QB (\$dummy [1007]), .D (nx41480), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41481 (.Y (nx41480), .A0 (ram_174__3), .A1 (nx65822), .S0 (
             nx63448)) ;
    oai21 ix58828 (.Y (nx58827), .A0 (nx10196), .A1 (nx10118), .B0 (nx65226)) ;
    nand04 ix10197 (.Y (nx10196), .A0 (nx58830), .A1 (nx58838), .A2 (nx58846), .A3 (
           nx58854)) ;
    aoi22 ix58831 (.Y (nx58830), .A0 (ram_176__3), .A1 (nx64506), .B0 (
          ram_177__3), .B1 (nx64544)) ;
    dffr reg_ram_176__3 (.Q (ram_176__3), .QB (\$dummy [1008]), .D (nx41460), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41461 (.Y (nx41460), .A0 (ram_176__3), .A1 (nx65822), .S0 (
             nx63434)) ;
    dffr reg_ram_177__3 (.Q (ram_177__3), .QB (\$dummy [1009]), .D (nx41450), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41451 (.Y (nx41450), .A0 (ram_177__3), .A1 (nx65822), .S0 (
             nx63424)) ;
    aoi22 ix58839 (.Y (nx58838), .A0 (ram_179__3), .A1 (nx64582), .B0 (
          ram_178__3), .B1 (nx64620)) ;
    dffr reg_ram_179__3 (.Q (ram_179__3), .QB (\$dummy [1010]), .D (nx41430), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41431 (.Y (nx41430), .A0 (ram_179__3), .A1 (nx65822), .S0 (
             nx63404)) ;
    dffr reg_ram_178__3 (.Q (ram_178__3), .QB (\$dummy [1011]), .D (nx41440), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41441 (.Y (nx41440), .A0 (ram_178__3), .A1 (nx65822), .S0 (
             nx63414)) ;
    aoi22 ix58847 (.Y (nx58846), .A0 (ram_180__3), .A1 (nx64658), .B0 (
          ram_181__3), .B1 (nx64696)) ;
    dffr reg_ram_180__3 (.Q (ram_180__3), .QB (\$dummy [1012]), .D (nx41420), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41421 (.Y (nx41420), .A0 (ram_180__3), .A1 (nx65822), .S0 (
             nx63394)) ;
    dffr reg_ram_181__3 (.Q (ram_181__3), .QB (\$dummy [1013]), .D (nx41410), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41411 (.Y (nx41410), .A0 (ram_181__3), .A1 (nx65824), .S0 (
             nx63384)) ;
    aoi22 ix58855 (.Y (nx58854), .A0 (ram_183__3), .A1 (nx64734), .B0 (
          ram_182__3), .B1 (nx64772)) ;
    dffr reg_ram_183__3 (.Q (ram_183__3), .QB (\$dummy [1014]), .D (nx41390), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41391 (.Y (nx41390), .A0 (ram_183__3), .A1 (nx65824), .S0 (
             nx63364)) ;
    dffr reg_ram_182__3 (.Q (ram_182__3), .QB (\$dummy [1015]), .D (nx41400), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41401 (.Y (nx41400), .A0 (ram_182__3), .A1 (nx65824), .S0 (
             nx63374)) ;
    nand04 ix10119 (.Y (nx10118), .A0 (nx58863), .A1 (nx58871), .A2 (nx58879), .A3 (
           nx58887)) ;
    aoi22 ix58864 (.Y (nx58863), .A0 (ram_184__3), .A1 (nx64810), .B0 (
          ram_185__3), .B1 (nx64848)) ;
    dffr reg_ram_184__3 (.Q (ram_184__3), .QB (\$dummy [1016]), .D (nx41380), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41381 (.Y (nx41380), .A0 (ram_184__3), .A1 (nx65824), .S0 (
             nx63354)) ;
    dffr reg_ram_185__3 (.Q (ram_185__3), .QB (\$dummy [1017]), .D (nx41370), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41371 (.Y (nx41370), .A0 (ram_185__3), .A1 (nx65824), .S0 (
             nx63344)) ;
    aoi22 ix58872 (.Y (nx58871), .A0 (ram_187__3), .A1 (nx64886), .B0 (
          ram_186__3), .B1 (nx64924)) ;
    dffr reg_ram_187__3 (.Q (ram_187__3), .QB (\$dummy [1018]), .D (nx41350), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41351 (.Y (nx41350), .A0 (ram_187__3), .A1 (nx65824), .S0 (
             nx63324)) ;
    dffr reg_ram_186__3 (.Q (ram_186__3), .QB (\$dummy [1019]), .D (nx41360), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41361 (.Y (nx41360), .A0 (ram_186__3), .A1 (nx65824), .S0 (
             nx63334)) ;
    aoi22 ix58880 (.Y (nx58879), .A0 (ram_188__3), .A1 (nx64962), .B0 (
          ram_189__3), .B1 (nx65000)) ;
    dffr reg_ram_188__3 (.Q (ram_188__3), .QB (\$dummy [1020]), .D (nx41340), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41341 (.Y (nx41340), .A0 (ram_188__3), .A1 (nx65826), .S0 (
             nx63314)) ;
    dffr reg_ram_189__3 (.Q (ram_189__3), .QB (\$dummy [1021]), .D (nx41330), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41331 (.Y (nx41330), .A0 (ram_189__3), .A1 (nx65826), .S0 (
             nx63304)) ;
    aoi22 ix58888 (.Y (nx58887), .A0 (ram_191__3), .A1 (nx65038), .B0 (
          ram_190__3), .B1 (nx65076)) ;
    dffr reg_ram_191__3 (.Q (ram_191__3), .QB (\$dummy [1022]), .D (nx41310), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41311 (.Y (nx41310), .A0 (ram_191__3), .A1 (nx65826), .S0 (
             nx63284)) ;
    dffr reg_ram_190__3 (.Q (ram_190__3), .QB (\$dummy [1023]), .D (nx41320), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix41321 (.Y (nx41320), .A0 (ram_190__3), .A1 (nx65826), .S0 (
             nx63294)) ;
    or04 ix15285 (.Y (dataout[4]), .A0 (nx15280), .A1 (nx14626), .A2 (nx13970), 
         .A3 (nx13316)) ;
    nand04 ix15281 (.Y (nx15280), .A0 (nx58897), .A1 (nx58965), .A2 (nx59033), .A3 (
           nx59101)) ;
    oai21 ix58898 (.Y (nx58897), .A0 (nx15270), .A1 (nx15192), .B0 (nx65096)) ;
    nand04 ix15271 (.Y (nx15270), .A0 (nx58900), .A1 (nx58908), .A2 (nx58916), .A3 (
           nx58924)) ;
    aoi22 ix58901 (.Y (nx58900), .A0 (ram_240__4), .A1 (nx64506), .B0 (
          ram_241__4), .B1 (nx64544)) ;
    dffr reg_ram_240__4 (.Q (ram_240__4), .QB (\$dummy [1024]), .D (nx46420), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46421 (.Y (nx46420), .A0 (ram_240__4), .A1 (nx65678), .S0 (
             nx64414)) ;
    dffr reg_ram_241__4 (.Q (ram_241__4), .QB (\$dummy [1025]), .D (nx46410), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46411 (.Y (nx46410), .A0 (ram_241__4), .A1 (nx65678), .S0 (
             nx64410)) ;
    aoi22 ix58909 (.Y (nx58908), .A0 (ram_243__4), .A1 (nx64582), .B0 (
          ram_242__4), .B1 (nx64620)) ;
    dffr reg_ram_243__4 (.Q (ram_243__4), .QB (\$dummy [1026]), .D (nx46390), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46391 (.Y (nx46390), .A0 (ram_243__4), .A1 (nx65678), .S0 (
             nx64402)) ;
    dffr reg_ram_242__4 (.Q (ram_242__4), .QB (\$dummy [1027]), .D (nx46400), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46401 (.Y (nx46400), .A0 (ram_242__4), .A1 (nx65678), .S0 (
             nx64406)) ;
    aoi22 ix58917 (.Y (nx58916), .A0 (ram_244__4), .A1 (nx64658), .B0 (
          ram_245__4), .B1 (nx64696)) ;
    dffr reg_ram_244__4 (.Q (ram_244__4), .QB (\$dummy [1028]), .D (nx46380), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46381 (.Y (nx46380), .A0 (ram_244__4), .A1 (nx65678), .S0 (
             nx64398)) ;
    dffr reg_ram_245__4 (.Q (ram_245__4), .QB (\$dummy [1029]), .D (nx46370), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46371 (.Y (nx46370), .A0 (ram_245__4), .A1 (nx65678), .S0 (
             nx64394)) ;
    aoi22 ix58925 (.Y (nx58924), .A0 (ram_247__4), .A1 (nx64734), .B0 (
          ram_246__4), .B1 (nx64772)) ;
    dffr reg_ram_247__4 (.Q (ram_247__4), .QB (\$dummy [1030]), .D (nx46350), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46351 (.Y (nx46350), .A0 (ram_247__4), .A1 (nx65678), .S0 (
             nx64386)) ;
    dffr reg_ram_246__4 (.Q (ram_246__4), .QB (\$dummy [1031]), .D (nx46360), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46361 (.Y (nx46360), .A0 (ram_246__4), .A1 (nx65680), .S0 (
             nx64390)) ;
    nand04 ix15193 (.Y (nx15192), .A0 (nx58933), .A1 (nx58941), .A2 (nx58949), .A3 (
           nx58957)) ;
    aoi22 ix58934 (.Y (nx58933), .A0 (ram_248__4), .A1 (nx64810), .B0 (
          ram_249__4), .B1 (nx64848)) ;
    dffr reg_ram_248__4 (.Q (ram_248__4), .QB (\$dummy [1032]), .D (nx46340), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46341 (.Y (nx46340), .A0 (ram_248__4), .A1 (nx65680), .S0 (
             nx64382)) ;
    dffr reg_ram_249__4 (.Q (ram_249__4), .QB (\$dummy [1033]), .D (nx46330), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46331 (.Y (nx46330), .A0 (ram_249__4), .A1 (nx65680), .S0 (
             nx64378)) ;
    aoi22 ix58942 (.Y (nx58941), .A0 (ram_251__4), .A1 (nx64886), .B0 (
          ram_250__4), .B1 (nx64924)) ;
    dffr reg_ram_251__4 (.Q (ram_251__4), .QB (\$dummy [1034]), .D (nx46310), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46311 (.Y (nx46310), .A0 (ram_251__4), .A1 (nx65680), .S0 (
             nx64370)) ;
    dffr reg_ram_250__4 (.Q (ram_250__4), .QB (\$dummy [1035]), .D (nx46320), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46321 (.Y (nx46320), .A0 (ram_250__4), .A1 (nx65680), .S0 (
             nx64374)) ;
    aoi22 ix58950 (.Y (nx58949), .A0 (ram_252__4), .A1 (nx64962), .B0 (
          ram_253__4), .B1 (nx65000)) ;
    dffr reg_ram_252__4 (.Q (ram_252__4), .QB (\$dummy [1036]), .D (nx46300), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46301 (.Y (nx46300), .A0 (ram_252__4), .A1 (nx65680), .S0 (
             nx64366)) ;
    dffr reg_ram_253__4 (.Q (ram_253__4), .QB (\$dummy [1037]), .D (nx46290), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46291 (.Y (nx46290), .A0 (ram_253__4), .A1 (nx65680), .S0 (
             nx64362)) ;
    aoi22 ix58958 (.Y (nx58957), .A0 (ram_255__4), .A1 (nx65038), .B0 (
          ram_254__4), .B1 (nx65076)) ;
    dffr reg_ram_255__4 (.Q (ram_255__4), .QB (\$dummy [1038]), .D (nx46270), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46271 (.Y (nx46270), .A0 (ram_255__4), .A1 (nx65682), .S0 (
             nx64354)) ;
    dffr reg_ram_254__4 (.Q (ram_254__4), .QB (\$dummy [1039]), .D (nx46280), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46281 (.Y (nx46280), .A0 (ram_254__4), .A1 (nx65682), .S0 (
             nx64358)) ;
    oai21 ix58966 (.Y (nx58965), .A0 (nx15108), .A1 (nx15030), .B0 (nx65100)) ;
    nand04 ix15109 (.Y (nx15108), .A0 (nx58968), .A1 (nx58976), .A2 (nx58984), .A3 (
           nx58992)) ;
    aoi22 ix58969 (.Y (nx58968), .A0 (ram_224__4), .A1 (nx64506), .B0 (
          ram_225__4), .B1 (nx64544)) ;
    dffr reg_ram_224__4 (.Q (ram_224__4), .QB (\$dummy [1040]), .D (nx46260), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46261 (.Y (nx46260), .A0 (ram_224__4), .A1 (nx65682), .S0 (
             nx64344)) ;
    dffr reg_ram_225__4 (.Q (ram_225__4), .QB (\$dummy [1041]), .D (nx46250), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46251 (.Y (nx46250), .A0 (ram_225__4), .A1 (nx65682), .S0 (
             nx64340)) ;
    aoi22 ix58977 (.Y (nx58976), .A0 (ram_227__4), .A1 (nx64582), .B0 (
          ram_226__4), .B1 (nx64620)) ;
    dffr reg_ram_227__4 (.Q (ram_227__4), .QB (\$dummy [1042]), .D (nx46230), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46231 (.Y (nx46230), .A0 (ram_227__4), .A1 (nx65682), .S0 (
             nx64332)) ;
    dffr reg_ram_226__4 (.Q (ram_226__4), .QB (\$dummy [1043]), .D (nx46240), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46241 (.Y (nx46240), .A0 (ram_226__4), .A1 (nx65682), .S0 (
             nx64336)) ;
    aoi22 ix58985 (.Y (nx58984), .A0 (ram_228__4), .A1 (nx64658), .B0 (
          ram_229__4), .B1 (nx64696)) ;
    dffr reg_ram_228__4 (.Q (ram_228__4), .QB (\$dummy [1044]), .D (nx46220), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46221 (.Y (nx46220), .A0 (ram_228__4), .A1 (nx65682), .S0 (
             nx64328)) ;
    dffr reg_ram_229__4 (.Q (ram_229__4), .QB (\$dummy [1045]), .D (nx46210), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46211 (.Y (nx46210), .A0 (ram_229__4), .A1 (nx65684), .S0 (
             nx64324)) ;
    aoi22 ix58993 (.Y (nx58992), .A0 (ram_231__4), .A1 (nx64734), .B0 (
          ram_230__4), .B1 (nx64772)) ;
    dffr reg_ram_231__4 (.Q (ram_231__4), .QB (\$dummy [1046]), .D (nx46190), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46191 (.Y (nx46190), .A0 (ram_231__4), .A1 (nx65684), .S0 (
             nx64316)) ;
    dffr reg_ram_230__4 (.Q (ram_230__4), .QB (\$dummy [1047]), .D (nx46200), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46201 (.Y (nx46200), .A0 (ram_230__4), .A1 (nx65684), .S0 (
             nx64320)) ;
    nand04 ix15031 (.Y (nx15030), .A0 (nx59001), .A1 (nx59009), .A2 (nx59017), .A3 (
           nx59025)) ;
    aoi22 ix59002 (.Y (nx59001), .A0 (ram_232__4), .A1 (nx64810), .B0 (
          ram_233__4), .B1 (nx64848)) ;
    dffr reg_ram_232__4 (.Q (ram_232__4), .QB (\$dummy [1048]), .D (nx46180), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46181 (.Y (nx46180), .A0 (ram_232__4), .A1 (nx65684), .S0 (
             nx64312)) ;
    dffr reg_ram_233__4 (.Q (ram_233__4), .QB (\$dummy [1049]), .D (nx46170), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46171 (.Y (nx46170), .A0 (ram_233__4), .A1 (nx65684), .S0 (
             nx64308)) ;
    aoi22 ix59010 (.Y (nx59009), .A0 (ram_235__4), .A1 (nx64886), .B0 (
          ram_234__4), .B1 (nx64924)) ;
    dffr reg_ram_235__4 (.Q (ram_235__4), .QB (\$dummy [1050]), .D (nx46150), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46151 (.Y (nx46150), .A0 (ram_235__4), .A1 (nx65684), .S0 (
             nx64300)) ;
    dffr reg_ram_234__4 (.Q (ram_234__4), .QB (\$dummy [1051]), .D (nx46160), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46161 (.Y (nx46160), .A0 (ram_234__4), .A1 (nx65684), .S0 (
             nx64304)) ;
    aoi22 ix59018 (.Y (nx59017), .A0 (ram_236__4), .A1 (nx64962), .B0 (
          ram_237__4), .B1 (nx65000)) ;
    dffr reg_ram_236__4 (.Q (ram_236__4), .QB (\$dummy [1052]), .D (nx46140), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46141 (.Y (nx46140), .A0 (ram_236__4), .A1 (nx65686), .S0 (
             nx64296)) ;
    dffr reg_ram_237__4 (.Q (ram_237__4), .QB (\$dummy [1053]), .D (nx46130), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46131 (.Y (nx46130), .A0 (ram_237__4), .A1 (nx65686), .S0 (
             nx64292)) ;
    aoi22 ix59026 (.Y (nx59025), .A0 (ram_239__4), .A1 (nx65038), .B0 (
          ram_238__4), .B1 (nx65076)) ;
    dffr reg_ram_239__4 (.Q (ram_239__4), .QB (\$dummy [1054]), .D (nx46110), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46111 (.Y (nx46110), .A0 (ram_239__4), .A1 (nx65686), .S0 (
             nx64284)) ;
    dffr reg_ram_238__4 (.Q (ram_238__4), .QB (\$dummy [1055]), .D (nx46120), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46121 (.Y (nx46120), .A0 (ram_238__4), .A1 (nx65686), .S0 (
             nx64288)) ;
    oai21 ix59034 (.Y (nx59033), .A0 (nx14944), .A1 (nx14866), .B0 (nx65104)) ;
    nand04 ix14945 (.Y (nx14944), .A0 (nx59036), .A1 (nx59044), .A2 (nx59052), .A3 (
           nx59060)) ;
    aoi22 ix59037 (.Y (nx59036), .A0 (ram_208__4), .A1 (nx64506), .B0 (
          ram_209__4), .B1 (nx64544)) ;
    dffr reg_ram_208__4 (.Q (ram_208__4), .QB (\$dummy [1056]), .D (nx46100), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46101 (.Y (nx46100), .A0 (ram_208__4), .A1 (nx65686), .S0 (
             nx64274)) ;
    dffr reg_ram_209__4 (.Q (ram_209__4), .QB (\$dummy [1057]), .D (nx46090), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46091 (.Y (nx46090), .A0 (ram_209__4), .A1 (nx65686), .S0 (
             nx64270)) ;
    aoi22 ix59045 (.Y (nx59044), .A0 (ram_211__4), .A1 (nx64582), .B0 (
          ram_210__4), .B1 (nx64620)) ;
    dffr reg_ram_211__4 (.Q (ram_211__4), .QB (\$dummy [1058]), .D (nx46070), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46071 (.Y (nx46070), .A0 (ram_211__4), .A1 (nx65686), .S0 (
             nx64262)) ;
    dffr reg_ram_210__4 (.Q (ram_210__4), .QB (\$dummy [1059]), .D (nx46080), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46081 (.Y (nx46080), .A0 (ram_210__4), .A1 (nx65688), .S0 (
             nx64266)) ;
    aoi22 ix59053 (.Y (nx59052), .A0 (ram_212__4), .A1 (nx64658), .B0 (
          ram_213__4), .B1 (nx64696)) ;
    dffr reg_ram_212__4 (.Q (ram_212__4), .QB (\$dummy [1060]), .D (nx46060), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46061 (.Y (nx46060), .A0 (ram_212__4), .A1 (nx65688), .S0 (
             nx64258)) ;
    dffr reg_ram_213__4 (.Q (ram_213__4), .QB (\$dummy [1061]), .D (nx46050), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46051 (.Y (nx46050), .A0 (ram_213__4), .A1 (nx65688), .S0 (
             nx64254)) ;
    aoi22 ix59061 (.Y (nx59060), .A0 (ram_215__4), .A1 (nx64734), .B0 (
          ram_214__4), .B1 (nx64772)) ;
    dffr reg_ram_215__4 (.Q (ram_215__4), .QB (\$dummy [1062]), .D (nx46030), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46031 (.Y (nx46030), .A0 (ram_215__4), .A1 (nx65688), .S0 (
             nx64246)) ;
    dffr reg_ram_214__4 (.Q (ram_214__4), .QB (\$dummy [1063]), .D (nx46040), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46041 (.Y (nx46040), .A0 (ram_214__4), .A1 (nx65688), .S0 (
             nx64250)) ;
    nand04 ix14867 (.Y (nx14866), .A0 (nx59069), .A1 (nx59077), .A2 (nx59085), .A3 (
           nx59093)) ;
    aoi22 ix59070 (.Y (nx59069), .A0 (ram_216__4), .A1 (nx64810), .B0 (
          ram_217__4), .B1 (nx64848)) ;
    dffr reg_ram_216__4 (.Q (ram_216__4), .QB (\$dummy [1064]), .D (nx46020), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46021 (.Y (nx46020), .A0 (ram_216__4), .A1 (nx65688), .S0 (
             nx64242)) ;
    dffr reg_ram_217__4 (.Q (ram_217__4), .QB (\$dummy [1065]), .D (nx46010), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46011 (.Y (nx46010), .A0 (ram_217__4), .A1 (nx65688), .S0 (
             nx64238)) ;
    aoi22 ix59078 (.Y (nx59077), .A0 (ram_219__4), .A1 (nx64886), .B0 (
          ram_218__4), .B1 (nx64924)) ;
    dffr reg_ram_219__4 (.Q (ram_219__4), .QB (\$dummy [1066]), .D (nx45990), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45991 (.Y (nx45990), .A0 (ram_219__4), .A1 (nx65690), .S0 (
             nx64230)) ;
    dffr reg_ram_218__4 (.Q (ram_218__4), .QB (\$dummy [1067]), .D (nx46000), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46001 (.Y (nx46000), .A0 (ram_218__4), .A1 (nx65690), .S0 (
             nx64234)) ;
    aoi22 ix59086 (.Y (nx59085), .A0 (ram_220__4), .A1 (nx64962), .B0 (
          ram_221__4), .B1 (nx65000)) ;
    dffr reg_ram_220__4 (.Q (ram_220__4), .QB (\$dummy [1068]), .D (nx45980), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45981 (.Y (nx45980), .A0 (ram_220__4), .A1 (nx65690), .S0 (
             nx64226)) ;
    dffr reg_ram_221__4 (.Q (ram_221__4), .QB (\$dummy [1069]), .D (nx45970), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45971 (.Y (nx45970), .A0 (ram_221__4), .A1 (nx65690), .S0 (
             nx64222)) ;
    aoi22 ix59094 (.Y (nx59093), .A0 (ram_223__4), .A1 (nx65038), .B0 (
          ram_222__4), .B1 (nx65076)) ;
    dffr reg_ram_223__4 (.Q (ram_223__4), .QB (\$dummy [1070]), .D (nx45950), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45951 (.Y (nx45950), .A0 (ram_223__4), .A1 (nx65690), .S0 (
             nx64214)) ;
    dffr reg_ram_222__4 (.Q (ram_222__4), .QB (\$dummy [1071]), .D (nx45960), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45961 (.Y (nx45960), .A0 (ram_222__4), .A1 (nx65690), .S0 (
             nx64218)) ;
    oai21 ix59102 (.Y (nx59101), .A0 (nx14782), .A1 (nx14704), .B0 (nx65108)) ;
    nand04 ix14783 (.Y (nx14782), .A0 (nx59104), .A1 (nx59112), .A2 (nx59120), .A3 (
           nx59128)) ;
    aoi22 ix59105 (.Y (nx59104), .A0 (ram_192__4), .A1 (nx64506), .B0 (
          ram_193__4), .B1 (nx64544)) ;
    dffr reg_ram_192__4 (.Q (ram_192__4), .QB (\$dummy [1072]), .D (nx45940), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45941 (.Y (nx45940), .A0 (ram_192__4), .A1 (nx65690), .S0 (
             nx64204)) ;
    dffr reg_ram_193__4 (.Q (ram_193__4), .QB (\$dummy [1073]), .D (nx45930), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45931 (.Y (nx45930), .A0 (ram_193__4), .A1 (nx65692), .S0 (
             nx64200)) ;
    aoi22 ix59113 (.Y (nx59112), .A0 (ram_195__4), .A1 (nx64582), .B0 (
          ram_194__4), .B1 (nx64620)) ;
    dffr reg_ram_195__4 (.Q (ram_195__4), .QB (\$dummy [1074]), .D (nx45910), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45911 (.Y (nx45910), .A0 (ram_195__4), .A1 (nx65692), .S0 (
             nx64192)) ;
    dffr reg_ram_194__4 (.Q (ram_194__4), .QB (\$dummy [1075]), .D (nx45920), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45921 (.Y (nx45920), .A0 (ram_194__4), .A1 (nx65692), .S0 (
             nx64196)) ;
    aoi22 ix59121 (.Y (nx59120), .A0 (ram_196__4), .A1 (nx64658), .B0 (
          ram_197__4), .B1 (nx64696)) ;
    dffr reg_ram_196__4 (.Q (ram_196__4), .QB (\$dummy [1076]), .D (nx45900), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45901 (.Y (nx45900), .A0 (ram_196__4), .A1 (nx65692), .S0 (
             nx64188)) ;
    dffr reg_ram_197__4 (.Q (ram_197__4), .QB (\$dummy [1077]), .D (nx45890), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45891 (.Y (nx45890), .A0 (ram_197__4), .A1 (nx65692), .S0 (
             nx64184)) ;
    aoi22 ix59129 (.Y (nx59128), .A0 (ram_199__4), .A1 (nx64734), .B0 (
          ram_198__4), .B1 (nx64772)) ;
    dffr reg_ram_199__4 (.Q (ram_199__4), .QB (\$dummy [1078]), .D (nx45870), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45871 (.Y (nx45870), .A0 (ram_199__4), .A1 (nx65692), .S0 (
             nx64176)) ;
    dffr reg_ram_198__4 (.Q (ram_198__4), .QB (\$dummy [1079]), .D (nx45880), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45881 (.Y (nx45880), .A0 (ram_198__4), .A1 (nx65692), .S0 (
             nx64180)) ;
    nand04 ix14705 (.Y (nx14704), .A0 (nx59137), .A1 (nx59145), .A2 (nx59153), .A3 (
           nx59161)) ;
    aoi22 ix59138 (.Y (nx59137), .A0 (ram_200__4), .A1 (nx64810), .B0 (
          ram_201__4), .B1 (nx64848)) ;
    dffr reg_ram_200__4 (.Q (ram_200__4), .QB (\$dummy [1080]), .D (nx45860), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45861 (.Y (nx45860), .A0 (ram_200__4), .A1 (nx65694), .S0 (
             nx64172)) ;
    dffr reg_ram_201__4 (.Q (ram_201__4), .QB (\$dummy [1081]), .D (nx45850), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45851 (.Y (nx45850), .A0 (ram_201__4), .A1 (nx65694), .S0 (
             nx64168)) ;
    aoi22 ix59146 (.Y (nx59145), .A0 (ram_203__4), .A1 (nx64886), .B0 (
          ram_202__4), .B1 (nx64924)) ;
    dffr reg_ram_203__4 (.Q (ram_203__4), .QB (\$dummy [1082]), .D (nx45830), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45831 (.Y (nx45830), .A0 (ram_203__4), .A1 (nx65694), .S0 (
             nx64160)) ;
    dffr reg_ram_202__4 (.Q (ram_202__4), .QB (\$dummy [1083]), .D (nx45840), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45841 (.Y (nx45840), .A0 (ram_202__4), .A1 (nx65694), .S0 (
             nx64164)) ;
    aoi22 ix59154 (.Y (nx59153), .A0 (ram_204__4), .A1 (nx64962), .B0 (
          ram_205__4), .B1 (nx65000)) ;
    dffr reg_ram_204__4 (.Q (ram_204__4), .QB (\$dummy [1084]), .D (nx45820), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45821 (.Y (nx45820), .A0 (ram_204__4), .A1 (nx65694), .S0 (
             nx64156)) ;
    dffr reg_ram_205__4 (.Q (ram_205__4), .QB (\$dummy [1085]), .D (nx45810), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45811 (.Y (nx45810), .A0 (ram_205__4), .A1 (nx65694), .S0 (
             nx64152)) ;
    aoi22 ix59162 (.Y (nx59161), .A0 (ram_207__4), .A1 (nx65038), .B0 (
          ram_206__4), .B1 (nx65076)) ;
    dffr reg_ram_207__4 (.Q (ram_207__4), .QB (\$dummy [1086]), .D (nx45790), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45791 (.Y (nx45790), .A0 (ram_207__4), .A1 (nx65694), .S0 (
             nx64144)) ;
    dffr reg_ram_206__4 (.Q (ram_206__4), .QB (\$dummy [1087]), .D (nx45800), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45801 (.Y (nx45800), .A0 (ram_206__4), .A1 (nx65696), .S0 (
             nx64148)) ;
    nand04 ix14627 (.Y (nx14626), .A0 (nx59170), .A1 (nx59238), .A2 (nx59306), .A3 (
           nx59374)) ;
    oai21 ix59171 (.Y (nx59170), .A0 (nx14616), .A1 (nx14538), .B0 (nx65112)) ;
    nand04 ix14617 (.Y (nx14616), .A0 (nx59173), .A1 (nx59181), .A2 (nx59189), .A3 (
           nx59197)) ;
    aoi22 ix59174 (.Y (nx59173), .A0 (ram_80__4), .A1 (nx64506), .B0 (ram_81__4)
          , .B1 (nx64544)) ;
    dffr reg_ram_80__4 (.Q (ram_80__4), .QB (\$dummy [1088]), .D (nx45780), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45781 (.Y (nx45780), .A0 (ram_80__4), .A1 (nx65696), .S0 (nx64134
             )) ;
    dffr reg_ram_81__4 (.Q (ram_81__4), .QB (\$dummy [1089]), .D (nx45770), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45771 (.Y (nx45770), .A0 (ram_81__4), .A1 (nx65696), .S0 (nx64130
             )) ;
    aoi22 ix59182 (.Y (nx59181), .A0 (ram_83__4), .A1 (nx64582), .B0 (ram_82__4)
          , .B1 (nx64620)) ;
    dffr reg_ram_83__4 (.Q (ram_83__4), .QB (\$dummy [1090]), .D (nx45750), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45751 (.Y (nx45750), .A0 (ram_83__4), .A1 (nx65696), .S0 (nx64122
             )) ;
    dffr reg_ram_82__4 (.Q (ram_82__4), .QB (\$dummy [1091]), .D (nx45760), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45761 (.Y (nx45760), .A0 (ram_82__4), .A1 (nx65696), .S0 (nx64126
             )) ;
    aoi22 ix59190 (.Y (nx59189), .A0 (ram_84__4), .A1 (nx64658), .B0 (ram_85__4)
          , .B1 (nx64696)) ;
    dffr reg_ram_84__4 (.Q (ram_84__4), .QB (\$dummy [1092]), .D (nx45740), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45741 (.Y (nx45740), .A0 (ram_84__4), .A1 (nx65696), .S0 (nx64118
             )) ;
    dffr reg_ram_85__4 (.Q (ram_85__4), .QB (\$dummy [1093]), .D (nx45730), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45731 (.Y (nx45730), .A0 (ram_85__4), .A1 (nx65696), .S0 (nx64114
             )) ;
    aoi22 ix59198 (.Y (nx59197), .A0 (ram_87__4), .A1 (nx64734), .B0 (ram_86__4)
          , .B1 (nx64772)) ;
    dffr reg_ram_87__4 (.Q (ram_87__4), .QB (\$dummy [1094]), .D (nx45710), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45711 (.Y (nx45710), .A0 (ram_87__4), .A1 (nx65698), .S0 (nx64106
             )) ;
    dffr reg_ram_86__4 (.Q (ram_86__4), .QB (\$dummy [1095]), .D (nx45720), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45721 (.Y (nx45720), .A0 (ram_86__4), .A1 (nx65698), .S0 (nx64110
             )) ;
    nand04 ix14539 (.Y (nx14538), .A0 (nx59206), .A1 (nx59214), .A2 (nx59222), .A3 (
           nx59230)) ;
    aoi22 ix59207 (.Y (nx59206), .A0 (ram_88__4), .A1 (nx64810), .B0 (ram_89__4)
          , .B1 (nx64848)) ;
    dffr reg_ram_88__4 (.Q (ram_88__4), .QB (\$dummy [1096]), .D (nx45700), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45701 (.Y (nx45700), .A0 (ram_88__4), .A1 (nx65698), .S0 (nx64102
             )) ;
    dffr reg_ram_89__4 (.Q (ram_89__4), .QB (\$dummy [1097]), .D (nx45690), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45691 (.Y (nx45690), .A0 (ram_89__4), .A1 (nx65698), .S0 (nx64098
             )) ;
    aoi22 ix59215 (.Y (nx59214), .A0 (ram_91__4), .A1 (nx64886), .B0 (ram_90__4)
          , .B1 (nx64924)) ;
    dffr reg_ram_91__4 (.Q (ram_91__4), .QB (\$dummy [1098]), .D (nx45670), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45671 (.Y (nx45670), .A0 (ram_91__4), .A1 (nx65698), .S0 (nx64090
             )) ;
    dffr reg_ram_90__4 (.Q (ram_90__4), .QB (\$dummy [1099]), .D (nx45680), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45681 (.Y (nx45680), .A0 (ram_90__4), .A1 (nx65698), .S0 (nx64094
             )) ;
    aoi22 ix59223 (.Y (nx59222), .A0 (ram_92__4), .A1 (nx64962), .B0 (ram_93__4)
          , .B1 (nx65000)) ;
    dffr reg_ram_92__4 (.Q (ram_92__4), .QB (\$dummy [1100]), .D (nx45660), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45661 (.Y (nx45660), .A0 (ram_92__4), .A1 (nx65698), .S0 (nx64086
             )) ;
    dffr reg_ram_93__4 (.Q (ram_93__4), .QB (\$dummy [1101]), .D (nx45650), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45651 (.Y (nx45650), .A0 (ram_93__4), .A1 (nx65700), .S0 (nx64082
             )) ;
    aoi22 ix59231 (.Y (nx59230), .A0 (ram_95__4), .A1 (nx65038), .B0 (ram_94__4)
          , .B1 (nx65076)) ;
    dffr reg_ram_95__4 (.Q (ram_95__4), .QB (\$dummy [1102]), .D (nx45630), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45631 (.Y (nx45630), .A0 (ram_95__4), .A1 (nx65700), .S0 (nx64074
             )) ;
    dffr reg_ram_94__4 (.Q (ram_94__4), .QB (\$dummy [1103]), .D (nx45640), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45641 (.Y (nx45640), .A0 (ram_94__4), .A1 (nx65700), .S0 (nx64078
             )) ;
    oai21 ix59239 (.Y (nx59238), .A0 (nx14454), .A1 (nx14376), .B0 (nx65116)) ;
    nand04 ix14455 (.Y (nx14454), .A0 (nx59241), .A1 (nx59249), .A2 (nx59257), .A3 (
           nx59265)) ;
    aoi22 ix59242 (.Y (nx59241), .A0 (ram_64__4), .A1 (nx64508), .B0 (ram_65__4)
          , .B1 (nx64546)) ;
    dffr reg_ram_64__4 (.Q (ram_64__4), .QB (\$dummy [1104]), .D (nx45620), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45621 (.Y (nx45620), .A0 (ram_64__4), .A1 (nx65700), .S0 (nx64064
             )) ;
    dffr reg_ram_65__4 (.Q (ram_65__4), .QB (\$dummy [1105]), .D (nx45610), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45611 (.Y (nx45610), .A0 (ram_65__4), .A1 (nx65700), .S0 (nx64060
             )) ;
    aoi22 ix59250 (.Y (nx59249), .A0 (ram_67__4), .A1 (nx64584), .B0 (ram_66__4)
          , .B1 (nx64622)) ;
    dffr reg_ram_67__4 (.Q (ram_67__4), .QB (\$dummy [1106]), .D (nx45590), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45591 (.Y (nx45590), .A0 (ram_67__4), .A1 (nx65700), .S0 (nx64052
             )) ;
    dffr reg_ram_66__4 (.Q (ram_66__4), .QB (\$dummy [1107]), .D (nx45600), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45601 (.Y (nx45600), .A0 (ram_66__4), .A1 (nx65700), .S0 (nx64056
             )) ;
    aoi22 ix59258 (.Y (nx59257), .A0 (ram_68__4), .A1 (nx64660), .B0 (ram_69__4)
          , .B1 (nx64698)) ;
    dffr reg_ram_68__4 (.Q (ram_68__4), .QB (\$dummy [1108]), .D (nx45580), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45581 (.Y (nx45580), .A0 (ram_68__4), .A1 (nx65702), .S0 (nx64048
             )) ;
    dffr reg_ram_69__4 (.Q (ram_69__4), .QB (\$dummy [1109]), .D (nx45570), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45571 (.Y (nx45570), .A0 (ram_69__4), .A1 (nx65702), .S0 (nx64044
             )) ;
    aoi22 ix59266 (.Y (nx59265), .A0 (ram_71__4), .A1 (nx64736), .B0 (ram_70__4)
          , .B1 (nx64774)) ;
    dffr reg_ram_71__4 (.Q (ram_71__4), .QB (\$dummy [1110]), .D (nx45550), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45551 (.Y (nx45550), .A0 (ram_71__4), .A1 (nx65702), .S0 (nx64036
             )) ;
    dffr reg_ram_70__4 (.Q (ram_70__4), .QB (\$dummy [1111]), .D (nx45560), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45561 (.Y (nx45560), .A0 (ram_70__4), .A1 (nx65702), .S0 (nx64040
             )) ;
    nand04 ix14377 (.Y (nx14376), .A0 (nx59274), .A1 (nx59282), .A2 (nx59290), .A3 (
           nx59298)) ;
    aoi22 ix59275 (.Y (nx59274), .A0 (ram_72__4), .A1 (nx64812), .B0 (ram_73__4)
          , .B1 (nx64850)) ;
    dffr reg_ram_72__4 (.Q (ram_72__4), .QB (\$dummy [1112]), .D (nx45540), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45541 (.Y (nx45540), .A0 (ram_72__4), .A1 (nx65702), .S0 (nx64032
             )) ;
    dffr reg_ram_73__4 (.Q (ram_73__4), .QB (\$dummy [1113]), .D (nx45530), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45531 (.Y (nx45530), .A0 (ram_73__4), .A1 (nx65702), .S0 (nx64028
             )) ;
    aoi22 ix59283 (.Y (nx59282), .A0 (ram_75__4), .A1 (nx64888), .B0 (ram_74__4)
          , .B1 (nx64926)) ;
    dffr reg_ram_75__4 (.Q (ram_75__4), .QB (\$dummy [1114]), .D (nx45510), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45511 (.Y (nx45510), .A0 (ram_75__4), .A1 (nx65702), .S0 (nx64020
             )) ;
    dffr reg_ram_74__4 (.Q (ram_74__4), .QB (\$dummy [1115]), .D (nx45520), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45521 (.Y (nx45520), .A0 (ram_74__4), .A1 (nx65704), .S0 (nx64024
             )) ;
    aoi22 ix59291 (.Y (nx59290), .A0 (ram_76__4), .A1 (nx64964), .B0 (ram_77__4)
          , .B1 (nx65002)) ;
    dffr reg_ram_76__4 (.Q (ram_76__4), .QB (\$dummy [1116]), .D (nx45500), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45501 (.Y (nx45500), .A0 (ram_76__4), .A1 (nx65704), .S0 (nx64016
             )) ;
    dffr reg_ram_77__4 (.Q (ram_77__4), .QB (\$dummy [1117]), .D (nx45490), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45491 (.Y (nx45490), .A0 (ram_77__4), .A1 (nx65704), .S0 (nx64012
             )) ;
    aoi22 ix59299 (.Y (nx59298), .A0 (ram_79__4), .A1 (nx65040), .B0 (ram_78__4)
          , .B1 (nx65078)) ;
    dffr reg_ram_79__4 (.Q (ram_79__4), .QB (\$dummy [1118]), .D (nx45470), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45471 (.Y (nx45470), .A0 (ram_79__4), .A1 (nx65704), .S0 (nx64004
             )) ;
    dffr reg_ram_78__4 (.Q (ram_78__4), .QB (\$dummy [1119]), .D (nx45480), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45481 (.Y (nx45480), .A0 (ram_78__4), .A1 (nx65704), .S0 (nx64008
             )) ;
    oai21 ix59307 (.Y (nx59306), .A0 (nx14290), .A1 (nx14212), .B0 (nx65120)) ;
    nand04 ix14291 (.Y (nx14290), .A0 (nx59309), .A1 (nx59317), .A2 (nx59325), .A3 (
           nx59333)) ;
    aoi22 ix59310 (.Y (nx59309), .A0 (ram_48__4), .A1 (nx64508), .B0 (ram_49__4)
          , .B1 (nx64546)) ;
    dffr reg_ram_48__4 (.Q (ram_48__4), .QB (\$dummy [1120]), .D (nx45460), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45461 (.Y (nx45460), .A0 (ram_48__4), .A1 (nx65704), .S0 (nx63994
             )) ;
    dffr reg_ram_49__4 (.Q (ram_49__4), .QB (\$dummy [1121]), .D (nx45450), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45451 (.Y (nx45450), .A0 (ram_49__4), .A1 (nx65704), .S0 (nx63990
             )) ;
    aoi22 ix59318 (.Y (nx59317), .A0 (ram_51__4), .A1 (nx64584), .B0 (ram_50__4)
          , .B1 (nx64622)) ;
    dffr reg_ram_51__4 (.Q (ram_51__4), .QB (\$dummy [1122]), .D (nx45430), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45431 (.Y (nx45430), .A0 (ram_51__4), .A1 (nx65706), .S0 (nx63982
             )) ;
    dffr reg_ram_50__4 (.Q (ram_50__4), .QB (\$dummy [1123]), .D (nx45440), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45441 (.Y (nx45440), .A0 (ram_50__4), .A1 (nx65706), .S0 (nx63986
             )) ;
    aoi22 ix59326 (.Y (nx59325), .A0 (ram_52__4), .A1 (nx64660), .B0 (ram_53__4)
          , .B1 (nx64698)) ;
    dffr reg_ram_52__4 (.Q (ram_52__4), .QB (\$dummy [1124]), .D (nx45420), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45421 (.Y (nx45420), .A0 (ram_52__4), .A1 (nx65706), .S0 (nx63978
             )) ;
    dffr reg_ram_53__4 (.Q (ram_53__4), .QB (\$dummy [1125]), .D (nx45410), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45411 (.Y (nx45410), .A0 (ram_53__4), .A1 (nx65706), .S0 (nx63974
             )) ;
    aoi22 ix59334 (.Y (nx59333), .A0 (ram_55__4), .A1 (nx64736), .B0 (ram_54__4)
          , .B1 (nx64774)) ;
    dffr reg_ram_55__4 (.Q (ram_55__4), .QB (\$dummy [1126]), .D (nx45390), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45391 (.Y (nx45390), .A0 (ram_55__4), .A1 (nx65706), .S0 (nx63966
             )) ;
    dffr reg_ram_54__4 (.Q (ram_54__4), .QB (\$dummy [1127]), .D (nx45400), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45401 (.Y (nx45400), .A0 (ram_54__4), .A1 (nx65706), .S0 (nx63970
             )) ;
    nand04 ix14213 (.Y (nx14212), .A0 (nx59342), .A1 (nx59350), .A2 (nx59358), .A3 (
           nx59366)) ;
    aoi22 ix59343 (.Y (nx59342), .A0 (ram_56__4), .A1 (nx64812), .B0 (ram_57__4)
          , .B1 (nx64850)) ;
    dffr reg_ram_56__4 (.Q (ram_56__4), .QB (\$dummy [1128]), .D (nx45380), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45381 (.Y (nx45380), .A0 (ram_56__4), .A1 (nx65706), .S0 (nx63962
             )) ;
    dffr reg_ram_57__4 (.Q (ram_57__4), .QB (\$dummy [1129]), .D (nx45370), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45371 (.Y (nx45370), .A0 (ram_57__4), .A1 (nx65708), .S0 (nx63958
             )) ;
    aoi22 ix59351 (.Y (nx59350), .A0 (ram_59__4), .A1 (nx64888), .B0 (ram_58__4)
          , .B1 (nx64926)) ;
    dffr reg_ram_59__4 (.Q (ram_59__4), .QB (\$dummy [1130]), .D (nx45350), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45351 (.Y (nx45350), .A0 (ram_59__4), .A1 (nx65708), .S0 (nx63950
             )) ;
    dffr reg_ram_58__4 (.Q (ram_58__4), .QB (\$dummy [1131]), .D (nx45360), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45361 (.Y (nx45360), .A0 (ram_58__4), .A1 (nx65708), .S0 (nx63954
             )) ;
    aoi22 ix59359 (.Y (nx59358), .A0 (ram_60__4), .A1 (nx64964), .B0 (ram_61__4)
          , .B1 (nx65002)) ;
    dffr reg_ram_60__4 (.Q (ram_60__4), .QB (\$dummy [1132]), .D (nx45340), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45341 (.Y (nx45340), .A0 (ram_60__4), .A1 (nx65708), .S0 (nx63946
             )) ;
    dffr reg_ram_61__4 (.Q (ram_61__4), .QB (\$dummy [1133]), .D (nx45330), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45331 (.Y (nx45330), .A0 (ram_61__4), .A1 (nx65708), .S0 (nx63942
             )) ;
    aoi22 ix59367 (.Y (nx59366), .A0 (ram_63__4), .A1 (nx65040), .B0 (ram_62__4)
          , .B1 (nx65078)) ;
    dffr reg_ram_63__4 (.Q (ram_63__4), .QB (\$dummy [1134]), .D (nx45310), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45311 (.Y (nx45310), .A0 (ram_63__4), .A1 (nx65708), .S0 (nx63934
             )) ;
    dffr reg_ram_62__4 (.Q (ram_62__4), .QB (\$dummy [1135]), .D (nx45320), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45321 (.Y (nx45320), .A0 (ram_62__4), .A1 (nx65708), .S0 (nx63938
             )) ;
    oai21 ix59375 (.Y (nx59374), .A0 (nx14128), .A1 (nx14050), .B0 (nx65124)) ;
    nand04 ix14129 (.Y (nx14128), .A0 (nx59377), .A1 (nx59385), .A2 (nx59393), .A3 (
           nx59401)) ;
    aoi22 ix59378 (.Y (nx59377), .A0 (ram_32__4), .A1 (nx64508), .B0 (ram_33__4)
          , .B1 (nx64546)) ;
    dffr reg_ram_32__4 (.Q (ram_32__4), .QB (\$dummy [1136]), .D (nx45300), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45301 (.Y (nx45300), .A0 (ram_32__4), .A1 (nx65710), .S0 (nx63924
             )) ;
    dffr reg_ram_33__4 (.Q (ram_33__4), .QB (\$dummy [1137]), .D (nx45290), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45291 (.Y (nx45290), .A0 (ram_33__4), .A1 (nx65710), .S0 (nx63920
             )) ;
    aoi22 ix59386 (.Y (nx59385), .A0 (ram_35__4), .A1 (nx64584), .B0 (ram_34__4)
          , .B1 (nx64622)) ;
    dffr reg_ram_35__4 (.Q (ram_35__4), .QB (\$dummy [1138]), .D (nx45270), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45271 (.Y (nx45270), .A0 (ram_35__4), .A1 (nx65710), .S0 (nx63912
             )) ;
    dffr reg_ram_34__4 (.Q (ram_34__4), .QB (\$dummy [1139]), .D (nx45280), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45281 (.Y (nx45280), .A0 (ram_34__4), .A1 (nx65710), .S0 (nx63916
             )) ;
    aoi22 ix59394 (.Y (nx59393), .A0 (ram_36__4), .A1 (nx64660), .B0 (ram_37__4)
          , .B1 (nx64698)) ;
    dffr reg_ram_36__4 (.Q (ram_36__4), .QB (\$dummy [1140]), .D (nx45260), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45261 (.Y (nx45260), .A0 (ram_36__4), .A1 (nx65710), .S0 (nx63908
             )) ;
    dffr reg_ram_37__4 (.Q (ram_37__4), .QB (\$dummy [1141]), .D (nx45250), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45251 (.Y (nx45250), .A0 (ram_37__4), .A1 (nx65710), .S0 (nx63904
             )) ;
    aoi22 ix59402 (.Y (nx59401), .A0 (ram_39__4), .A1 (nx64736), .B0 (ram_38__4)
          , .B1 (nx64774)) ;
    dffr reg_ram_39__4 (.Q (ram_39__4), .QB (\$dummy [1142]), .D (nx45230), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45231 (.Y (nx45230), .A0 (ram_39__4), .A1 (nx65710), .S0 (nx63896
             )) ;
    dffr reg_ram_38__4 (.Q (ram_38__4), .QB (\$dummy [1143]), .D (nx45240), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45241 (.Y (nx45240), .A0 (ram_38__4), .A1 (nx65712), .S0 (nx63900
             )) ;
    nand04 ix14051 (.Y (nx14050), .A0 (nx59410), .A1 (nx59418), .A2 (nx59426), .A3 (
           nx59434)) ;
    aoi22 ix59411 (.Y (nx59410), .A0 (ram_40__4), .A1 (nx64812), .B0 (ram_41__4)
          , .B1 (nx64850)) ;
    dffr reg_ram_40__4 (.Q (ram_40__4), .QB (\$dummy [1144]), .D (nx45220), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45221 (.Y (nx45220), .A0 (ram_40__4), .A1 (nx65712), .S0 (nx63892
             )) ;
    dffr reg_ram_41__4 (.Q (ram_41__4), .QB (\$dummy [1145]), .D (nx45210), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45211 (.Y (nx45210), .A0 (ram_41__4), .A1 (nx65712), .S0 (nx63888
             )) ;
    aoi22 ix59419 (.Y (nx59418), .A0 (ram_43__4), .A1 (nx64888), .B0 (ram_42__4)
          , .B1 (nx64926)) ;
    dffr reg_ram_43__4 (.Q (ram_43__4), .QB (\$dummy [1146]), .D (nx45190), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45191 (.Y (nx45190), .A0 (ram_43__4), .A1 (nx65712), .S0 (nx63880
             )) ;
    dffr reg_ram_42__4 (.Q (ram_42__4), .QB (\$dummy [1147]), .D (nx45200), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45201 (.Y (nx45200), .A0 (ram_42__4), .A1 (nx65712), .S0 (nx63884
             )) ;
    aoi22 ix59427 (.Y (nx59426), .A0 (ram_44__4), .A1 (nx64964), .B0 (ram_45__4)
          , .B1 (nx65002)) ;
    dffr reg_ram_44__4 (.Q (ram_44__4), .QB (\$dummy [1148]), .D (nx45180), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45181 (.Y (nx45180), .A0 (ram_44__4), .A1 (nx65712), .S0 (nx63876
             )) ;
    dffr reg_ram_45__4 (.Q (ram_45__4), .QB (\$dummy [1149]), .D (nx45170), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45171 (.Y (nx45170), .A0 (ram_45__4), .A1 (nx65712), .S0 (nx63872
             )) ;
    aoi22 ix59435 (.Y (nx59434), .A0 (ram_47__4), .A1 (nx65040), .B0 (ram_46__4)
          , .B1 (nx65078)) ;
    dffr reg_ram_47__4 (.Q (ram_47__4), .QB (\$dummy [1150]), .D (nx45150), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45151 (.Y (nx45150), .A0 (ram_47__4), .A1 (nx65714), .S0 (nx63864
             )) ;
    dffr reg_ram_46__4 (.Q (ram_46__4), .QB (\$dummy [1151]), .D (nx45160), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45161 (.Y (nx45160), .A0 (ram_46__4), .A1 (nx65714), .S0 (nx63868
             )) ;
    nand04 ix13971 (.Y (nx13970), .A0 (nx59443), .A1 (nx59511), .A2 (nx59579), .A3 (
           nx59647)) ;
    oai21 ix59444 (.Y (nx59443), .A0 (nx13960), .A1 (nx13882), .B0 (nx65128)) ;
    nand04 ix13961 (.Y (nx13960), .A0 (nx59446), .A1 (nx59454), .A2 (nx59462), .A3 (
           nx59470)) ;
    aoi22 ix59447 (.Y (nx59446), .A0 (ram_16__4), .A1 (nx64508), .B0 (ram_17__4)
          , .B1 (nx64546)) ;
    dffr reg_ram_16__4 (.Q (ram_16__4), .QB (\$dummy [1152]), .D (nx45140), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45141 (.Y (nx45140), .A0 (ram_16__4), .A1 (nx65714), .S0 (nx63854
             )) ;
    dffr reg_ram_17__4 (.Q (ram_17__4), .QB (\$dummy [1153]), .D (nx45130), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45131 (.Y (nx45130), .A0 (ram_17__4), .A1 (nx65714), .S0 (nx63850
             )) ;
    aoi22 ix59455 (.Y (nx59454), .A0 (ram_19__4), .A1 (nx64584), .B0 (ram_18__4)
          , .B1 (nx64622)) ;
    dffr reg_ram_19__4 (.Q (ram_19__4), .QB (\$dummy [1154]), .D (nx45110), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45111 (.Y (nx45110), .A0 (ram_19__4), .A1 (nx65714), .S0 (nx63842
             )) ;
    dffr reg_ram_18__4 (.Q (ram_18__4), .QB (\$dummy [1155]), .D (nx45120), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45121 (.Y (nx45120), .A0 (ram_18__4), .A1 (nx65714), .S0 (nx63846
             )) ;
    aoi22 ix59463 (.Y (nx59462), .A0 (ram_20__4), .A1 (nx64660), .B0 (ram_21__4)
          , .B1 (nx64698)) ;
    dffr reg_ram_20__4 (.Q (ram_20__4), .QB (\$dummy [1156]), .D (nx45100), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45101 (.Y (nx45100), .A0 (ram_20__4), .A1 (nx65714), .S0 (nx63838
             )) ;
    dffr reg_ram_21__4 (.Q (ram_21__4), .QB (\$dummy [1157]), .D (nx45090), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45091 (.Y (nx45090), .A0 (ram_21__4), .A1 (nx65716), .S0 (nx63834
             )) ;
    aoi22 ix59471 (.Y (nx59470), .A0 (ram_23__4), .A1 (nx64736), .B0 (ram_22__4)
          , .B1 (nx64774)) ;
    dffr reg_ram_23__4 (.Q (ram_23__4), .QB (\$dummy [1158]), .D (nx45070), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45071 (.Y (nx45070), .A0 (ram_23__4), .A1 (nx65716), .S0 (nx63826
             )) ;
    dffr reg_ram_22__4 (.Q (ram_22__4), .QB (\$dummy [1159]), .D (nx45080), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45081 (.Y (nx45080), .A0 (ram_22__4), .A1 (nx65716), .S0 (nx63830
             )) ;
    nand04 ix13883 (.Y (nx13882), .A0 (nx59479), .A1 (nx59487), .A2 (nx59495), .A3 (
           nx59503)) ;
    aoi22 ix59480 (.Y (nx59479), .A0 (ram_24__4), .A1 (nx64812), .B0 (ram_25__4)
          , .B1 (nx64850)) ;
    dffr reg_ram_24__4 (.Q (ram_24__4), .QB (\$dummy [1160]), .D (nx45060), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45061 (.Y (nx45060), .A0 (ram_24__4), .A1 (nx65716), .S0 (nx63822
             )) ;
    dffr reg_ram_25__4 (.Q (ram_25__4), .QB (\$dummy [1161]), .D (nx45050), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45051 (.Y (nx45050), .A0 (ram_25__4), .A1 (nx65716), .S0 (nx63818
             )) ;
    aoi22 ix59488 (.Y (nx59487), .A0 (ram_27__4), .A1 (nx64888), .B0 (ram_26__4)
          , .B1 (nx64926)) ;
    dffr reg_ram_27__4 (.Q (ram_27__4), .QB (\$dummy [1162]), .D (nx45030), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45031 (.Y (nx45030), .A0 (ram_27__4), .A1 (nx65716), .S0 (nx63810
             )) ;
    dffr reg_ram_26__4 (.Q (ram_26__4), .QB (\$dummy [1163]), .D (nx45040), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45041 (.Y (nx45040), .A0 (ram_26__4), .A1 (nx65716), .S0 (nx63814
             )) ;
    aoi22 ix59496 (.Y (nx59495), .A0 (ram_28__4), .A1 (nx64964), .B0 (ram_29__4)
          , .B1 (nx65002)) ;
    dffr reg_ram_28__4 (.Q (ram_28__4), .QB (\$dummy [1164]), .D (nx45020), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45021 (.Y (nx45020), .A0 (ram_28__4), .A1 (nx65718), .S0 (nx63806
             )) ;
    dffr reg_ram_29__4 (.Q (ram_29__4), .QB (\$dummy [1165]), .D (nx45010), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45011 (.Y (nx45010), .A0 (ram_29__4), .A1 (nx65718), .S0 (nx63802
             )) ;
    aoi22 ix59504 (.Y (nx59503), .A0 (ram_31__4), .A1 (nx65040), .B0 (ram_30__4)
          , .B1 (nx65078)) ;
    dffr reg_ram_31__4 (.Q (ram_31__4), .QB (\$dummy [1166]), .D (nx44990), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44991 (.Y (nx44990), .A0 (ram_31__4), .A1 (nx65718), .S0 (nx63794
             )) ;
    dffr reg_ram_30__4 (.Q (ram_30__4), .QB (\$dummy [1167]), .D (nx45000), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix45001 (.Y (nx45000), .A0 (ram_30__4), .A1 (nx65718), .S0 (nx63798
             )) ;
    oai21 ix59512 (.Y (nx59511), .A0 (nx13798), .A1 (nx13720), .B0 (nx65142)) ;
    nand04 ix13799 (.Y (nx13798), .A0 (nx59514), .A1 (nx59522), .A2 (nx59530), .A3 (
           nx59538)) ;
    aoi22 ix59515 (.Y (nx59514), .A0 (ram_0__4), .A1 (nx64508), .B0 (ram_1__4), 
          .B1 (nx64546)) ;
    dffr reg_ram_0__4 (.Q (ram_0__4), .QB (\$dummy [1168]), .D (nx44980), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44981 (.Y (nx44980), .A0 (nx65718), .A1 (ram_0__4), .S0 (nx65132)
             ) ;
    dffr reg_ram_1__4 (.Q (ram_1__4), .QB (\$dummy [1169]), .D (nx44970), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44971 (.Y (nx44970), .A0 (nx65718), .A1 (ram_1__4), .S0 (nx65146)
             ) ;
    aoi22 ix59523 (.Y (nx59522), .A0 (ram_3__4), .A1 (nx64584), .B0 (ram_2__4), 
          .B1 (nx64622)) ;
    dffr reg_ram_3__4 (.Q (ram_3__4), .QB (\$dummy [1170]), .D (nx44950), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44951 (.Y (nx44950), .A0 (nx65718), .A1 (ram_3__4), .S0 (nx65150)
             ) ;
    dffr reg_ram_2__4 (.Q (ram_2__4), .QB (\$dummy [1171]), .D (nx44960), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44961 (.Y (nx44960), .A0 (nx65720), .A1 (ram_2__4), .S0 (nx65154)
             ) ;
    aoi22 ix59531 (.Y (nx59530), .A0 (ram_4__4), .A1 (nx64660), .B0 (ram_5__4), 
          .B1 (nx64698)) ;
    dffr reg_ram_4__4 (.Q (ram_4__4), .QB (\$dummy [1172]), .D (nx44940), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44941 (.Y (nx44940), .A0 (nx65720), .A1 (ram_4__4), .S0 (nx65158)
             ) ;
    dffr reg_ram_5__4 (.Q (ram_5__4), .QB (\$dummy [1173]), .D (nx44930), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44931 (.Y (nx44930), .A0 (nx65720), .A1 (ram_5__4), .S0 (nx65162)
             ) ;
    aoi22 ix59539 (.Y (nx59538), .A0 (ram_7__4), .A1 (nx64736), .B0 (ram_6__4), 
          .B1 (nx64774)) ;
    dffr reg_ram_7__4 (.Q (ram_7__4), .QB (\$dummy [1174]), .D (nx44910), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44911 (.Y (nx44910), .A0 (nx65720), .A1 (ram_7__4), .S0 (nx65166)
             ) ;
    dffr reg_ram_6__4 (.Q (ram_6__4), .QB (\$dummy [1175]), .D (nx44920), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44921 (.Y (nx44920), .A0 (nx65720), .A1 (ram_6__4), .S0 (nx65170)
             ) ;
    nand04 ix13721 (.Y (nx13720), .A0 (nx59547), .A1 (nx59555), .A2 (nx59563), .A3 (
           nx59571)) ;
    aoi22 ix59548 (.Y (nx59547), .A0 (ram_8__4), .A1 (nx64812), .B0 (ram_9__4), 
          .B1 (nx64850)) ;
    dffr reg_ram_8__4 (.Q (ram_8__4), .QB (\$dummy [1176]), .D (nx44900), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44901 (.Y (nx44900), .A0 (nx65720), .A1 (ram_8__4), .S0 (nx65174)
             ) ;
    dffr reg_ram_9__4 (.Q (ram_9__4), .QB (\$dummy [1177]), .D (nx44890), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44891 (.Y (nx44890), .A0 (nx65720), .A1 (ram_9__4), .S0 (nx65178)
             ) ;
    aoi22 ix59556 (.Y (nx59555), .A0 (ram_11__4), .A1 (nx64888), .B0 (ram_10__4)
          , .B1 (nx64926)) ;
    dffr reg_ram_11__4 (.Q (ram_11__4), .QB (\$dummy [1178]), .D (nx44870), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44871 (.Y (nx44870), .A0 (nx65722), .A1 (ram_11__4), .S0 (nx65182
             )) ;
    dffr reg_ram_10__4 (.Q (ram_10__4), .QB (\$dummy [1179]), .D (nx44880), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44881 (.Y (nx44880), .A0 (nx65722), .A1 (ram_10__4), .S0 (nx65186
             )) ;
    aoi22 ix59564 (.Y (nx59563), .A0 (ram_12__4), .A1 (nx64964), .B0 (ram_13__4)
          , .B1 (nx65002)) ;
    dffr reg_ram_12__4 (.Q (ram_12__4), .QB (\$dummy [1180]), .D (nx44860), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44861 (.Y (nx44860), .A0 (nx65722), .A1 (ram_12__4), .S0 (nx65190
             )) ;
    dffr reg_ram_13__4 (.Q (ram_13__4), .QB (\$dummy [1181]), .D (nx44850), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44851 (.Y (nx44850), .A0 (nx65722), .A1 (ram_13__4), .S0 (nx65194
             )) ;
    aoi22 ix59572 (.Y (nx59571), .A0 (ram_15__4), .A1 (nx65040), .B0 (ram_14__4)
          , .B1 (nx65078)) ;
    dffr reg_ram_15__4 (.Q (ram_15__4), .QB (\$dummy [1182]), .D (nx44830), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44831 (.Y (nx44830), .A0 (nx65722), .A1 (ram_15__4), .S0 (nx65198
             )) ;
    dffr reg_ram_14__4 (.Q (ram_14__4), .QB (\$dummy [1183]), .D (nx44840), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44841 (.Y (nx44840), .A0 (nx65722), .A1 (ram_14__4), .S0 (nx65202
             )) ;
    oai21 ix59580 (.Y (nx59579), .A0 (nx13634), .A1 (nx13556), .B0 (nx65206)) ;
    nand04 ix13635 (.Y (nx13634), .A0 (nx59582), .A1 (nx59590), .A2 (nx59598), .A3 (
           nx59606)) ;
    aoi22 ix59583 (.Y (nx59582), .A0 (ram_96__4), .A1 (nx64508), .B0 (ram_97__4)
          , .B1 (nx64546)) ;
    dffr reg_ram_96__4 (.Q (ram_96__4), .QB (\$dummy [1184]), .D (nx44820), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44821 (.Y (nx44820), .A0 (ram_96__4), .A1 (nx65722), .S0 (nx63784
             )) ;
    dffr reg_ram_97__4 (.Q (ram_97__4), .QB (\$dummy [1185]), .D (nx44810), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44811 (.Y (nx44810), .A0 (ram_97__4), .A1 (nx65724), .S0 (nx63780
             )) ;
    aoi22 ix59591 (.Y (nx59590), .A0 (ram_99__4), .A1 (nx64584), .B0 (ram_98__4)
          , .B1 (nx64622)) ;
    dffr reg_ram_99__4 (.Q (ram_99__4), .QB (\$dummy [1186]), .D (nx44790), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44791 (.Y (nx44790), .A0 (ram_99__4), .A1 (nx65724), .S0 (nx63772
             )) ;
    dffr reg_ram_98__4 (.Q (ram_98__4), .QB (\$dummy [1187]), .D (nx44800), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44801 (.Y (nx44800), .A0 (ram_98__4), .A1 (nx65724), .S0 (nx63776
             )) ;
    aoi22 ix59599 (.Y (nx59598), .A0 (ram_100__4), .A1 (nx64660), .B0 (
          ram_101__4), .B1 (nx64698)) ;
    dffr reg_ram_100__4 (.Q (ram_100__4), .QB (\$dummy [1188]), .D (nx44780), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44781 (.Y (nx44780), .A0 (ram_100__4), .A1 (nx65724), .S0 (
             nx63768)) ;
    dffr reg_ram_101__4 (.Q (ram_101__4), .QB (\$dummy [1189]), .D (nx44770), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44771 (.Y (nx44770), .A0 (ram_101__4), .A1 (nx65724), .S0 (
             nx63764)) ;
    aoi22 ix59607 (.Y (nx59606), .A0 (ram_103__4), .A1 (nx64736), .B0 (
          ram_102__4), .B1 (nx64774)) ;
    dffr reg_ram_103__4 (.Q (ram_103__4), .QB (\$dummy [1190]), .D (nx44750), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44751 (.Y (nx44750), .A0 (ram_103__4), .A1 (nx65724), .S0 (
             nx63756)) ;
    dffr reg_ram_102__4 (.Q (ram_102__4), .QB (\$dummy [1191]), .D (nx44760), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44761 (.Y (nx44760), .A0 (ram_102__4), .A1 (nx65724), .S0 (
             nx63760)) ;
    nand04 ix13557 (.Y (nx13556), .A0 (nx59615), .A1 (nx59623), .A2 (nx59631), .A3 (
           nx59639)) ;
    aoi22 ix59616 (.Y (nx59615), .A0 (ram_104__4), .A1 (nx64812), .B0 (
          ram_105__4), .B1 (nx64850)) ;
    dffr reg_ram_104__4 (.Q (ram_104__4), .QB (\$dummy [1192]), .D (nx44740), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44741 (.Y (nx44740), .A0 (ram_104__4), .A1 (nx65726), .S0 (
             nx63752)) ;
    dffr reg_ram_105__4 (.Q (ram_105__4), .QB (\$dummy [1193]), .D (nx44730), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44731 (.Y (nx44730), .A0 (ram_105__4), .A1 (nx65726), .S0 (
             nx63748)) ;
    aoi22 ix59624 (.Y (nx59623), .A0 (ram_107__4), .A1 (nx64888), .B0 (
          ram_106__4), .B1 (nx64926)) ;
    dffr reg_ram_107__4 (.Q (ram_107__4), .QB (\$dummy [1194]), .D (nx44710), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44711 (.Y (nx44710), .A0 (ram_107__4), .A1 (nx65726), .S0 (
             nx63740)) ;
    dffr reg_ram_106__4 (.Q (ram_106__4), .QB (\$dummy [1195]), .D (nx44720), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44721 (.Y (nx44720), .A0 (ram_106__4), .A1 (nx65726), .S0 (
             nx63744)) ;
    aoi22 ix59632 (.Y (nx59631), .A0 (ram_108__4), .A1 (nx64964), .B0 (
          ram_109__4), .B1 (nx65002)) ;
    dffr reg_ram_108__4 (.Q (ram_108__4), .QB (\$dummy [1196]), .D (nx44700), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44701 (.Y (nx44700), .A0 (ram_108__4), .A1 (nx65726), .S0 (
             nx63736)) ;
    dffr reg_ram_109__4 (.Q (ram_109__4), .QB (\$dummy [1197]), .D (nx44690), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44691 (.Y (nx44690), .A0 (ram_109__4), .A1 (nx65726), .S0 (
             nx63732)) ;
    aoi22 ix59640 (.Y (nx59639), .A0 (ram_111__4), .A1 (nx65040), .B0 (
          ram_110__4), .B1 (nx65078)) ;
    dffr reg_ram_111__4 (.Q (ram_111__4), .QB (\$dummy [1198]), .D (nx44670), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44671 (.Y (nx44670), .A0 (ram_111__4), .A1 (nx65726), .S0 (
             nx63724)) ;
    dffr reg_ram_110__4 (.Q (ram_110__4), .QB (\$dummy [1199]), .D (nx44680), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44681 (.Y (nx44680), .A0 (ram_110__4), .A1 (nx65728), .S0 (
             nx63728)) ;
    oai21 ix59648 (.Y (nx59647), .A0 (nx13472), .A1 (nx13394), .B0 (nx65210)) ;
    nand04 ix13473 (.Y (nx13472), .A0 (nx59650), .A1 (nx59658), .A2 (nx59666), .A3 (
           nx59674)) ;
    aoi22 ix59651 (.Y (nx59650), .A0 (ram_112__4), .A1 (nx64508), .B0 (
          ram_113__4), .B1 (nx64546)) ;
    dffr reg_ram_112__4 (.Q (ram_112__4), .QB (\$dummy [1200]), .D (nx44660), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44661 (.Y (nx44660), .A0 (ram_112__4), .A1 (nx65728), .S0 (
             nx63714)) ;
    dffr reg_ram_113__4 (.Q (ram_113__4), .QB (\$dummy [1201]), .D (nx44650), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44651 (.Y (nx44650), .A0 (ram_113__4), .A1 (nx65728), .S0 (
             nx63710)) ;
    aoi22 ix59659 (.Y (nx59658), .A0 (ram_115__4), .A1 (nx64584), .B0 (
          ram_114__4), .B1 (nx64622)) ;
    dffr reg_ram_115__4 (.Q (ram_115__4), .QB (\$dummy [1202]), .D (nx44630), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44631 (.Y (nx44630), .A0 (ram_115__4), .A1 (nx65728), .S0 (
             nx63702)) ;
    dffr reg_ram_114__4 (.Q (ram_114__4), .QB (\$dummy [1203]), .D (nx44640), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44641 (.Y (nx44640), .A0 (ram_114__4), .A1 (nx65728), .S0 (
             nx63706)) ;
    aoi22 ix59667 (.Y (nx59666), .A0 (ram_116__4), .A1 (nx64660), .B0 (
          ram_117__4), .B1 (nx64698)) ;
    dffr reg_ram_116__4 (.Q (ram_116__4), .QB (\$dummy [1204]), .D (nx44620), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44621 (.Y (nx44620), .A0 (ram_116__4), .A1 (nx65728), .S0 (
             nx63698)) ;
    dffr reg_ram_117__4 (.Q (ram_117__4), .QB (\$dummy [1205]), .D (nx44610), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44611 (.Y (nx44610), .A0 (ram_117__4), .A1 (nx65728), .S0 (
             nx63694)) ;
    aoi22 ix59675 (.Y (nx59674), .A0 (ram_119__4), .A1 (nx64736), .B0 (
          ram_118__4), .B1 (nx64774)) ;
    dffr reg_ram_119__4 (.Q (ram_119__4), .QB (\$dummy [1206]), .D (nx44590), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44591 (.Y (nx44590), .A0 (ram_119__4), .A1 (nx65730), .S0 (
             nx63686)) ;
    dffr reg_ram_118__4 (.Q (ram_118__4), .QB (\$dummy [1207]), .D (nx44600), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44601 (.Y (nx44600), .A0 (ram_118__4), .A1 (nx65730), .S0 (
             nx63690)) ;
    nand04 ix13395 (.Y (nx13394), .A0 (nx59683), .A1 (nx59691), .A2 (nx59699), .A3 (
           nx59707)) ;
    aoi22 ix59684 (.Y (nx59683), .A0 (ram_120__4), .A1 (nx64812), .B0 (
          ram_121__4), .B1 (nx64850)) ;
    dffr reg_ram_120__4 (.Q (ram_120__4), .QB (\$dummy [1208]), .D (nx44580), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44581 (.Y (nx44580), .A0 (ram_120__4), .A1 (nx65730), .S0 (
             nx63682)) ;
    dffr reg_ram_121__4 (.Q (ram_121__4), .QB (\$dummy [1209]), .D (nx44570), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44571 (.Y (nx44570), .A0 (ram_121__4), .A1 (nx65730), .S0 (
             nx63678)) ;
    aoi22 ix59692 (.Y (nx59691), .A0 (ram_123__4), .A1 (nx64888), .B0 (
          ram_122__4), .B1 (nx64926)) ;
    dffr reg_ram_123__4 (.Q (ram_123__4), .QB (\$dummy [1210]), .D (nx44550), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44551 (.Y (nx44550), .A0 (ram_123__4), .A1 (nx65730), .S0 (
             nx63670)) ;
    dffr reg_ram_122__4 (.Q (ram_122__4), .QB (\$dummy [1211]), .D (nx44560), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44561 (.Y (nx44560), .A0 (ram_122__4), .A1 (nx65730), .S0 (
             nx63674)) ;
    aoi22 ix59700 (.Y (nx59699), .A0 (ram_124__4), .A1 (nx64964), .B0 (
          ram_125__4), .B1 (nx65002)) ;
    dffr reg_ram_124__4 (.Q (ram_124__4), .QB (\$dummy [1212]), .D (nx44540), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44541 (.Y (nx44540), .A0 (ram_124__4), .A1 (nx65730), .S0 (
             nx63666)) ;
    dffr reg_ram_125__4 (.Q (ram_125__4), .QB (\$dummy [1213]), .D (nx44530), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44531 (.Y (nx44530), .A0 (ram_125__4), .A1 (nx65732), .S0 (
             nx63662)) ;
    aoi22 ix59708 (.Y (nx59707), .A0 (ram_127__4), .A1 (nx65040), .B0 (
          ram_126__4), .B1 (nx65078)) ;
    dffr reg_ram_127__4 (.Q (ram_127__4), .QB (\$dummy [1214]), .D (nx44510), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44511 (.Y (nx44510), .A0 (ram_127__4), .A1 (nx65732), .S0 (
             nx63654)) ;
    dffr reg_ram_126__4 (.Q (ram_126__4), .QB (\$dummy [1215]), .D (nx44520), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44521 (.Y (nx44520), .A0 (ram_126__4), .A1 (nx65732), .S0 (
             nx63658)) ;
    nand04 ix13317 (.Y (nx13316), .A0 (nx59716), .A1 (nx59784), .A2 (nx59852), .A3 (
           nx59920)) ;
    oai21 ix59717 (.Y (nx59716), .A0 (nx13306), .A1 (nx13228), .B0 (nx65214)) ;
    nand04 ix13307 (.Y (nx13306), .A0 (nx59719), .A1 (nx59727), .A2 (nx59735), .A3 (
           nx59743)) ;
    aoi22 ix59720 (.Y (nx59719), .A0 (ram_128__4), .A1 (nx64510), .B0 (
          ram_129__4), .B1 (nx64548)) ;
    dffr reg_ram_128__4 (.Q (ram_128__4), .QB (\$dummy [1216]), .D (nx44500), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44501 (.Y (nx44500), .A0 (ram_128__4), .A1 (nx65732), .S0 (
             nx63644)) ;
    dffr reg_ram_129__4 (.Q (ram_129__4), .QB (\$dummy [1217]), .D (nx44490), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44491 (.Y (nx44490), .A0 (ram_129__4), .A1 (nx65732), .S0 (
             nx63640)) ;
    aoi22 ix59728 (.Y (nx59727), .A0 (ram_131__4), .A1 (nx64586), .B0 (
          ram_130__4), .B1 (nx64624)) ;
    dffr reg_ram_131__4 (.Q (ram_131__4), .QB (\$dummy [1218]), .D (nx44470), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44471 (.Y (nx44470), .A0 (ram_131__4), .A1 (nx65732), .S0 (
             nx63632)) ;
    dffr reg_ram_130__4 (.Q (ram_130__4), .QB (\$dummy [1219]), .D (nx44480), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44481 (.Y (nx44480), .A0 (ram_130__4), .A1 (nx65732), .S0 (
             nx63636)) ;
    aoi22 ix59736 (.Y (nx59735), .A0 (ram_132__4), .A1 (nx64662), .B0 (
          ram_133__4), .B1 (nx64700)) ;
    dffr reg_ram_132__4 (.Q (ram_132__4), .QB (\$dummy [1220]), .D (nx44460), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44461 (.Y (nx44460), .A0 (ram_132__4), .A1 (nx65734), .S0 (
             nx63628)) ;
    dffr reg_ram_133__4 (.Q (ram_133__4), .QB (\$dummy [1221]), .D (nx44450), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44451 (.Y (nx44450), .A0 (ram_133__4), .A1 (nx65734), .S0 (
             nx63624)) ;
    aoi22 ix59744 (.Y (nx59743), .A0 (ram_135__4), .A1 (nx64738), .B0 (
          ram_134__4), .B1 (nx64776)) ;
    dffr reg_ram_135__4 (.Q (ram_135__4), .QB (\$dummy [1222]), .D (nx44430), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44431 (.Y (nx44430), .A0 (ram_135__4), .A1 (nx65734), .S0 (
             nx63616)) ;
    dffr reg_ram_134__4 (.Q (ram_134__4), .QB (\$dummy [1223]), .D (nx44440), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44441 (.Y (nx44440), .A0 (ram_134__4), .A1 (nx65734), .S0 (
             nx63620)) ;
    nand04 ix13229 (.Y (nx13228), .A0 (nx59752), .A1 (nx59760), .A2 (nx59768), .A3 (
           nx59776)) ;
    aoi22 ix59753 (.Y (nx59752), .A0 (ram_136__4), .A1 (nx64814), .B0 (
          ram_137__4), .B1 (nx64852)) ;
    dffr reg_ram_136__4 (.Q (ram_136__4), .QB (\$dummy [1224]), .D (nx44420), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44421 (.Y (nx44420), .A0 (ram_136__4), .A1 (nx65734), .S0 (
             nx63612)) ;
    dffr reg_ram_137__4 (.Q (ram_137__4), .QB (\$dummy [1225]), .D (nx44410), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44411 (.Y (nx44410), .A0 (ram_137__4), .A1 (nx65734), .S0 (
             nx63608)) ;
    aoi22 ix59761 (.Y (nx59760), .A0 (ram_139__4), .A1 (nx64890), .B0 (
          ram_138__4), .B1 (nx64928)) ;
    dffr reg_ram_139__4 (.Q (ram_139__4), .QB (\$dummy [1226]), .D (nx44390), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44391 (.Y (nx44390), .A0 (ram_139__4), .A1 (nx65734), .S0 (
             nx63600)) ;
    dffr reg_ram_138__4 (.Q (ram_138__4), .QB (\$dummy [1227]), .D (nx44400), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44401 (.Y (nx44400), .A0 (ram_138__4), .A1 (nx65736), .S0 (
             nx63604)) ;
    aoi22 ix59769 (.Y (nx59768), .A0 (ram_140__4), .A1 (nx64966), .B0 (
          ram_141__4), .B1 (nx65004)) ;
    dffr reg_ram_140__4 (.Q (ram_140__4), .QB (\$dummy [1228]), .D (nx44380), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44381 (.Y (nx44380), .A0 (ram_140__4), .A1 (nx65736), .S0 (
             nx63596)) ;
    dffr reg_ram_141__4 (.Q (ram_141__4), .QB (\$dummy [1229]), .D (nx44370), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44371 (.Y (nx44370), .A0 (ram_141__4), .A1 (nx65736), .S0 (
             nx63592)) ;
    aoi22 ix59777 (.Y (nx59776), .A0 (ram_143__4), .A1 (nx65042), .B0 (
          ram_142__4), .B1 (nx65080)) ;
    dffr reg_ram_143__4 (.Q (ram_143__4), .QB (\$dummy [1230]), .D (nx44350), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44351 (.Y (nx44350), .A0 (ram_143__4), .A1 (nx65736), .S0 (
             nx63584)) ;
    dffr reg_ram_142__4 (.Q (ram_142__4), .QB (\$dummy [1231]), .D (nx44360), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44361 (.Y (nx44360), .A0 (ram_142__4), .A1 (nx65736), .S0 (
             nx63588)) ;
    oai21 ix59785 (.Y (nx59784), .A0 (nx13144), .A1 (nx13066), .B0 (nx65218)) ;
    nand04 ix13145 (.Y (nx13144), .A0 (nx59787), .A1 (nx59795), .A2 (nx59803), .A3 (
           nx59811)) ;
    aoi22 ix59788 (.Y (nx59787), .A0 (ram_144__4), .A1 (nx64510), .B0 (
          ram_145__4), .B1 (nx64548)) ;
    dffr reg_ram_144__4 (.Q (ram_144__4), .QB (\$dummy [1232]), .D (nx44340), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44341 (.Y (nx44340), .A0 (ram_144__4), .A1 (nx65736), .S0 (
             nx63574)) ;
    dffr reg_ram_145__4 (.Q (ram_145__4), .QB (\$dummy [1233]), .D (nx44330), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44331 (.Y (nx44330), .A0 (ram_145__4), .A1 (nx65736), .S0 (
             nx63570)) ;
    aoi22 ix59796 (.Y (nx59795), .A0 (ram_147__4), .A1 (nx64586), .B0 (
          ram_146__4), .B1 (nx64624)) ;
    dffr reg_ram_147__4 (.Q (ram_147__4), .QB (\$dummy [1234]), .D (nx44310), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44311 (.Y (nx44310), .A0 (ram_147__4), .A1 (nx65738), .S0 (
             nx63562)) ;
    dffr reg_ram_146__4 (.Q (ram_146__4), .QB (\$dummy [1235]), .D (nx44320), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44321 (.Y (nx44320), .A0 (ram_146__4), .A1 (nx65738), .S0 (
             nx63566)) ;
    aoi22 ix59804 (.Y (nx59803), .A0 (ram_148__4), .A1 (nx64662), .B0 (
          ram_149__4), .B1 (nx64700)) ;
    dffr reg_ram_148__4 (.Q (ram_148__4), .QB (\$dummy [1236]), .D (nx44300), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44301 (.Y (nx44300), .A0 (ram_148__4), .A1 (nx65738), .S0 (
             nx63558)) ;
    dffr reg_ram_149__4 (.Q (ram_149__4), .QB (\$dummy [1237]), .D (nx44290), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44291 (.Y (nx44290), .A0 (ram_149__4), .A1 (nx65738), .S0 (
             nx63554)) ;
    aoi22 ix59812 (.Y (nx59811), .A0 (ram_151__4), .A1 (nx64738), .B0 (
          ram_150__4), .B1 (nx64776)) ;
    dffr reg_ram_151__4 (.Q (ram_151__4), .QB (\$dummy [1238]), .D (nx44270), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44271 (.Y (nx44270), .A0 (ram_151__4), .A1 (nx65738), .S0 (
             nx63546)) ;
    dffr reg_ram_150__4 (.Q (ram_150__4), .QB (\$dummy [1239]), .D (nx44280), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44281 (.Y (nx44280), .A0 (ram_150__4), .A1 (nx65738), .S0 (
             nx63550)) ;
    nand04 ix13067 (.Y (nx13066), .A0 (nx59820), .A1 (nx59828), .A2 (nx59836), .A3 (
           nx59844)) ;
    aoi22 ix59821 (.Y (nx59820), .A0 (ram_152__4), .A1 (nx64814), .B0 (
          ram_153__4), .B1 (nx64852)) ;
    dffr reg_ram_152__4 (.Q (ram_152__4), .QB (\$dummy [1240]), .D (nx44260), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44261 (.Y (nx44260), .A0 (ram_152__4), .A1 (nx65738), .S0 (
             nx63542)) ;
    dffr reg_ram_153__4 (.Q (ram_153__4), .QB (\$dummy [1241]), .D (nx44250), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44251 (.Y (nx44250), .A0 (ram_153__4), .A1 (nx65740), .S0 (
             nx63538)) ;
    aoi22 ix59829 (.Y (nx59828), .A0 (ram_155__4), .A1 (nx64890), .B0 (
          ram_154__4), .B1 (nx64928)) ;
    dffr reg_ram_155__4 (.Q (ram_155__4), .QB (\$dummy [1242]), .D (nx44230), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44231 (.Y (nx44230), .A0 (ram_155__4), .A1 (nx65740), .S0 (
             nx63530)) ;
    dffr reg_ram_154__4 (.Q (ram_154__4), .QB (\$dummy [1243]), .D (nx44240), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44241 (.Y (nx44240), .A0 (ram_154__4), .A1 (nx65740), .S0 (
             nx63534)) ;
    aoi22 ix59837 (.Y (nx59836), .A0 (ram_156__4), .A1 (nx64966), .B0 (
          ram_157__4), .B1 (nx65004)) ;
    dffr reg_ram_156__4 (.Q (ram_156__4), .QB (\$dummy [1244]), .D (nx44220), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44221 (.Y (nx44220), .A0 (ram_156__4), .A1 (nx65740), .S0 (
             nx63526)) ;
    dffr reg_ram_157__4 (.Q (ram_157__4), .QB (\$dummy [1245]), .D (nx44210), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44211 (.Y (nx44210), .A0 (ram_157__4), .A1 (nx65740), .S0 (
             nx63522)) ;
    aoi22 ix59845 (.Y (nx59844), .A0 (ram_159__4), .A1 (nx65042), .B0 (
          ram_158__4), .B1 (nx65080)) ;
    dffr reg_ram_159__4 (.Q (ram_159__4), .QB (\$dummy [1246]), .D (nx44190), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44191 (.Y (nx44190), .A0 (ram_159__4), .A1 (nx65740), .S0 (
             nx63514)) ;
    dffr reg_ram_158__4 (.Q (ram_158__4), .QB (\$dummy [1247]), .D (nx44200), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44201 (.Y (nx44200), .A0 (ram_158__4), .A1 (nx65740), .S0 (
             nx63518)) ;
    oai21 ix59853 (.Y (nx59852), .A0 (nx12980), .A1 (nx12902), .B0 (nx65222)) ;
    nand04 ix12981 (.Y (nx12980), .A0 (nx59855), .A1 (nx59863), .A2 (nx59871), .A3 (
           nx59879)) ;
    aoi22 ix59856 (.Y (nx59855), .A0 (ram_160__4), .A1 (nx64510), .B0 (
          ram_161__4), .B1 (nx64548)) ;
    dffr reg_ram_160__4 (.Q (ram_160__4), .QB (\$dummy [1248]), .D (nx44180), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44181 (.Y (nx44180), .A0 (ram_160__4), .A1 (nx65742), .S0 (
             nx63504)) ;
    dffr reg_ram_161__4 (.Q (ram_161__4), .QB (\$dummy [1249]), .D (nx44170), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44171 (.Y (nx44170), .A0 (ram_161__4), .A1 (nx65742), .S0 (
             nx63500)) ;
    aoi22 ix59864 (.Y (nx59863), .A0 (ram_163__4), .A1 (nx64586), .B0 (
          ram_162__4), .B1 (nx64624)) ;
    dffr reg_ram_163__4 (.Q (ram_163__4), .QB (\$dummy [1250]), .D (nx44150), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44151 (.Y (nx44150), .A0 (ram_163__4), .A1 (nx65742), .S0 (
             nx63492)) ;
    dffr reg_ram_162__4 (.Q (ram_162__4), .QB (\$dummy [1251]), .D (nx44160), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44161 (.Y (nx44160), .A0 (ram_162__4), .A1 (nx65742), .S0 (
             nx63496)) ;
    aoi22 ix59872 (.Y (nx59871), .A0 (ram_164__4), .A1 (nx64662), .B0 (
          ram_165__4), .B1 (nx64700)) ;
    dffr reg_ram_164__4 (.Q (ram_164__4), .QB (\$dummy [1252]), .D (nx44140), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44141 (.Y (nx44140), .A0 (ram_164__4), .A1 (nx65742), .S0 (
             nx63488)) ;
    dffr reg_ram_165__4 (.Q (ram_165__4), .QB (\$dummy [1253]), .D (nx44130), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44131 (.Y (nx44130), .A0 (ram_165__4), .A1 (nx65742), .S0 (
             nx63484)) ;
    aoi22 ix59880 (.Y (nx59879), .A0 (ram_167__4), .A1 (nx64738), .B0 (
          ram_166__4), .B1 (nx64776)) ;
    dffr reg_ram_167__4 (.Q (ram_167__4), .QB (\$dummy [1254]), .D (nx44110), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44111 (.Y (nx44110), .A0 (ram_167__4), .A1 (nx65742), .S0 (
             nx63476)) ;
    dffr reg_ram_166__4 (.Q (ram_166__4), .QB (\$dummy [1255]), .D (nx44120), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44121 (.Y (nx44120), .A0 (ram_166__4), .A1 (nx65744), .S0 (
             nx63480)) ;
    nand04 ix12903 (.Y (nx12902), .A0 (nx59888), .A1 (nx59896), .A2 (nx59904), .A3 (
           nx59912)) ;
    aoi22 ix59889 (.Y (nx59888), .A0 (ram_168__4), .A1 (nx64814), .B0 (
          ram_169__4), .B1 (nx64852)) ;
    dffr reg_ram_168__4 (.Q (ram_168__4), .QB (\$dummy [1256]), .D (nx44100), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44101 (.Y (nx44100), .A0 (ram_168__4), .A1 (nx65744), .S0 (
             nx63472)) ;
    dffr reg_ram_169__4 (.Q (ram_169__4), .QB (\$dummy [1257]), .D (nx44090), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44091 (.Y (nx44090), .A0 (ram_169__4), .A1 (nx65744), .S0 (
             nx63468)) ;
    aoi22 ix59897 (.Y (nx59896), .A0 (ram_171__4), .A1 (nx64890), .B0 (
          ram_170__4), .B1 (nx64928)) ;
    dffr reg_ram_171__4 (.Q (ram_171__4), .QB (\$dummy [1258]), .D (nx44070), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44071 (.Y (nx44070), .A0 (ram_171__4), .A1 (nx65744), .S0 (
             nx63460)) ;
    dffr reg_ram_170__4 (.Q (ram_170__4), .QB (\$dummy [1259]), .D (nx44080), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44081 (.Y (nx44080), .A0 (ram_170__4), .A1 (nx65744), .S0 (
             nx63464)) ;
    aoi22 ix59905 (.Y (nx59904), .A0 (ram_172__4), .A1 (nx64966), .B0 (
          ram_173__4), .B1 (nx65004)) ;
    dffr reg_ram_172__4 (.Q (ram_172__4), .QB (\$dummy [1260]), .D (nx44060), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44061 (.Y (nx44060), .A0 (ram_172__4), .A1 (nx65744), .S0 (
             nx63456)) ;
    dffr reg_ram_173__4 (.Q (ram_173__4), .QB (\$dummy [1261]), .D (nx44050), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44051 (.Y (nx44050), .A0 (ram_173__4), .A1 (nx65744), .S0 (
             nx63452)) ;
    aoi22 ix59913 (.Y (nx59912), .A0 (ram_175__4), .A1 (nx65042), .B0 (
          ram_174__4), .B1 (nx65080)) ;
    dffr reg_ram_175__4 (.Q (ram_175__4), .QB (\$dummy [1262]), .D (nx44030), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44031 (.Y (nx44030), .A0 (ram_175__4), .A1 (nx65746), .S0 (
             nx63444)) ;
    dffr reg_ram_174__4 (.Q (ram_174__4), .QB (\$dummy [1263]), .D (nx44040), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44041 (.Y (nx44040), .A0 (ram_174__4), .A1 (nx65746), .S0 (
             nx63448)) ;
    oai21 ix59921 (.Y (nx59920), .A0 (nx12818), .A1 (nx12740), .B0 (nx65226)) ;
    nand04 ix12819 (.Y (nx12818), .A0 (nx59923), .A1 (nx59931), .A2 (nx59939), .A3 (
           nx59947)) ;
    aoi22 ix59924 (.Y (nx59923), .A0 (ram_176__4), .A1 (nx64510), .B0 (
          ram_177__4), .B1 (nx64548)) ;
    dffr reg_ram_176__4 (.Q (ram_176__4), .QB (\$dummy [1264]), .D (nx44020), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44021 (.Y (nx44020), .A0 (ram_176__4), .A1 (nx65746), .S0 (
             nx63434)) ;
    dffr reg_ram_177__4 (.Q (ram_177__4), .QB (\$dummy [1265]), .D (nx44010), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44011 (.Y (nx44010), .A0 (ram_177__4), .A1 (nx65746), .S0 (
             nx63424)) ;
    aoi22 ix59932 (.Y (nx59931), .A0 (ram_179__4), .A1 (nx64586), .B0 (
          ram_178__4), .B1 (nx64624)) ;
    dffr reg_ram_179__4 (.Q (ram_179__4), .QB (\$dummy [1266]), .D (nx43990), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43991 (.Y (nx43990), .A0 (ram_179__4), .A1 (nx65746), .S0 (
             nx63404)) ;
    dffr reg_ram_178__4 (.Q (ram_178__4), .QB (\$dummy [1267]), .D (nx44000), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix44001 (.Y (nx44000), .A0 (ram_178__4), .A1 (nx65746), .S0 (
             nx63414)) ;
    aoi22 ix59940 (.Y (nx59939), .A0 (ram_180__4), .A1 (nx64662), .B0 (
          ram_181__4), .B1 (nx64700)) ;
    dffr reg_ram_180__4 (.Q (ram_180__4), .QB (\$dummy [1268]), .D (nx43980), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43981 (.Y (nx43980), .A0 (ram_180__4), .A1 (nx65746), .S0 (
             nx63394)) ;
    dffr reg_ram_181__4 (.Q (ram_181__4), .QB (\$dummy [1269]), .D (nx43970), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43971 (.Y (nx43970), .A0 (ram_181__4), .A1 (nx65748), .S0 (
             nx63384)) ;
    aoi22 ix59948 (.Y (nx59947), .A0 (ram_183__4), .A1 (nx64738), .B0 (
          ram_182__4), .B1 (nx64776)) ;
    dffr reg_ram_183__4 (.Q (ram_183__4), .QB (\$dummy [1270]), .D (nx43950), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43951 (.Y (nx43950), .A0 (ram_183__4), .A1 (nx65748), .S0 (
             nx63364)) ;
    dffr reg_ram_182__4 (.Q (ram_182__4), .QB (\$dummy [1271]), .D (nx43960), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43961 (.Y (nx43960), .A0 (ram_182__4), .A1 (nx65748), .S0 (
             nx63374)) ;
    nand04 ix12741 (.Y (nx12740), .A0 (nx59956), .A1 (nx59964), .A2 (nx59972), .A3 (
           nx59980)) ;
    aoi22 ix59957 (.Y (nx59956), .A0 (ram_184__4), .A1 (nx64814), .B0 (
          ram_185__4), .B1 (nx64852)) ;
    dffr reg_ram_184__4 (.Q (ram_184__4), .QB (\$dummy [1272]), .D (nx43940), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43941 (.Y (nx43940), .A0 (ram_184__4), .A1 (nx65748), .S0 (
             nx63354)) ;
    dffr reg_ram_185__4 (.Q (ram_185__4), .QB (\$dummy [1273]), .D (nx43930), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43931 (.Y (nx43930), .A0 (ram_185__4), .A1 (nx65748), .S0 (
             nx63344)) ;
    aoi22 ix59965 (.Y (nx59964), .A0 (ram_187__4), .A1 (nx64890), .B0 (
          ram_186__4), .B1 (nx64928)) ;
    dffr reg_ram_187__4 (.Q (ram_187__4), .QB (\$dummy [1274]), .D (nx43910), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43911 (.Y (nx43910), .A0 (ram_187__4), .A1 (nx65748), .S0 (
             nx63324)) ;
    dffr reg_ram_186__4 (.Q (ram_186__4), .QB (\$dummy [1275]), .D (nx43920), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43921 (.Y (nx43920), .A0 (ram_186__4), .A1 (nx65748), .S0 (
             nx63334)) ;
    aoi22 ix59973 (.Y (nx59972), .A0 (ram_188__4), .A1 (nx64966), .B0 (
          ram_189__4), .B1 (nx65004)) ;
    dffr reg_ram_188__4 (.Q (ram_188__4), .QB (\$dummy [1276]), .D (nx43900), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43901 (.Y (nx43900), .A0 (ram_188__4), .A1 (nx65750), .S0 (
             nx63314)) ;
    dffr reg_ram_189__4 (.Q (ram_189__4), .QB (\$dummy [1277]), .D (nx43890), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43891 (.Y (nx43890), .A0 (ram_189__4), .A1 (nx65750), .S0 (
             nx63304)) ;
    aoi22 ix59981 (.Y (nx59980), .A0 (ram_191__4), .A1 (nx65042), .B0 (
          ram_190__4), .B1 (nx65080)) ;
    dffr reg_ram_191__4 (.Q (ram_191__4), .QB (\$dummy [1278]), .D (nx43870), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43871 (.Y (nx43870), .A0 (ram_191__4), .A1 (nx65750), .S0 (
             nx63284)) ;
    dffr reg_ram_190__4 (.Q (ram_190__4), .QB (\$dummy [1279]), .D (nx43880), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix43881 (.Y (nx43880), .A0 (ram_190__4), .A1 (nx65750), .S0 (
             nx63294)) ;
    or04 ix17907 (.Y (dataout[5]), .A0 (nx17902), .A1 (nx17248), .A2 (nx16592), 
         .A3 (nx15938)) ;
    nand04 ix17903 (.Y (nx17902), .A0 (nx59990), .A1 (nx60058), .A2 (nx60126), .A3 (
           nx60194)) ;
    oai21 ix59991 (.Y (nx59990), .A0 (nx17892), .A1 (nx17814), .B0 (nx65096)) ;
    nand04 ix17893 (.Y (nx17892), .A0 (nx59993), .A1 (nx60001), .A2 (nx60009), .A3 (
           nx60017)) ;
    aoi22 ix59994 (.Y (nx59993), .A0 (ram_240__5), .A1 (nx64510), .B0 (
          ram_241__5), .B1 (nx64548)) ;
    dffr reg_ram_240__5 (.Q (ram_240__5), .QB (\$dummy [1280]), .D (nx48980), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48981 (.Y (nx48980), .A0 (ram_240__5), .A1 (nx65602), .S0 (
             nx64414)) ;
    dffr reg_ram_241__5 (.Q (ram_241__5), .QB (\$dummy [1281]), .D (nx48970), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48971 (.Y (nx48970), .A0 (ram_241__5), .A1 (nx65602), .S0 (
             nx64410)) ;
    aoi22 ix60002 (.Y (nx60001), .A0 (ram_243__5), .A1 (nx64586), .B0 (
          ram_242__5), .B1 (nx64624)) ;
    dffr reg_ram_243__5 (.Q (ram_243__5), .QB (\$dummy [1282]), .D (nx48950), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48951 (.Y (nx48950), .A0 (ram_243__5), .A1 (nx65602), .S0 (
             nx64402)) ;
    dffr reg_ram_242__5 (.Q (ram_242__5), .QB (\$dummy [1283]), .D (nx48960), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48961 (.Y (nx48960), .A0 (ram_242__5), .A1 (nx65602), .S0 (
             nx64406)) ;
    aoi22 ix60010 (.Y (nx60009), .A0 (ram_244__5), .A1 (nx64662), .B0 (
          ram_245__5), .B1 (nx64700)) ;
    dffr reg_ram_244__5 (.Q (ram_244__5), .QB (\$dummy [1284]), .D (nx48940), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48941 (.Y (nx48940), .A0 (ram_244__5), .A1 (nx65602), .S0 (
             nx64398)) ;
    dffr reg_ram_245__5 (.Q (ram_245__5), .QB (\$dummy [1285]), .D (nx48930), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48931 (.Y (nx48930), .A0 (ram_245__5), .A1 (nx65602), .S0 (
             nx64394)) ;
    aoi22 ix60018 (.Y (nx60017), .A0 (ram_247__5), .A1 (nx64738), .B0 (
          ram_246__5), .B1 (nx64776)) ;
    dffr reg_ram_247__5 (.Q (ram_247__5), .QB (\$dummy [1286]), .D (nx48910), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48911 (.Y (nx48910), .A0 (ram_247__5), .A1 (nx65602), .S0 (
             nx64386)) ;
    dffr reg_ram_246__5 (.Q (ram_246__5), .QB (\$dummy [1287]), .D (nx48920), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48921 (.Y (nx48920), .A0 (ram_246__5), .A1 (nx65604), .S0 (
             nx64390)) ;
    nand04 ix17815 (.Y (nx17814), .A0 (nx60026), .A1 (nx60034), .A2 (nx60042), .A3 (
           nx60050)) ;
    aoi22 ix60027 (.Y (nx60026), .A0 (ram_248__5), .A1 (nx64814), .B0 (
          ram_249__5), .B1 (nx64852)) ;
    dffr reg_ram_248__5 (.Q (ram_248__5), .QB (\$dummy [1288]), .D (nx48900), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48901 (.Y (nx48900), .A0 (ram_248__5), .A1 (nx65604), .S0 (
             nx64382)) ;
    dffr reg_ram_249__5 (.Q (ram_249__5), .QB (\$dummy [1289]), .D (nx48890), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48891 (.Y (nx48890), .A0 (ram_249__5), .A1 (nx65604), .S0 (
             nx64378)) ;
    aoi22 ix60035 (.Y (nx60034), .A0 (ram_251__5), .A1 (nx64890), .B0 (
          ram_250__5), .B1 (nx64928)) ;
    dffr reg_ram_251__5 (.Q (ram_251__5), .QB (\$dummy [1290]), .D (nx48870), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48871 (.Y (nx48870), .A0 (ram_251__5), .A1 (nx65604), .S0 (
             nx64370)) ;
    dffr reg_ram_250__5 (.Q (ram_250__5), .QB (\$dummy [1291]), .D (nx48880), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48881 (.Y (nx48880), .A0 (ram_250__5), .A1 (nx65604), .S0 (
             nx64374)) ;
    aoi22 ix60043 (.Y (nx60042), .A0 (ram_252__5), .A1 (nx64966), .B0 (
          ram_253__5), .B1 (nx65004)) ;
    dffr reg_ram_252__5 (.Q (ram_252__5), .QB (\$dummy [1292]), .D (nx48860), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48861 (.Y (nx48860), .A0 (ram_252__5), .A1 (nx65604), .S0 (
             nx64366)) ;
    dffr reg_ram_253__5 (.Q (ram_253__5), .QB (\$dummy [1293]), .D (nx48850), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48851 (.Y (nx48850), .A0 (ram_253__5), .A1 (nx65604), .S0 (
             nx64362)) ;
    aoi22 ix60051 (.Y (nx60050), .A0 (ram_255__5), .A1 (nx65042), .B0 (
          ram_254__5), .B1 (nx65080)) ;
    dffr reg_ram_255__5 (.Q (ram_255__5), .QB (\$dummy [1294]), .D (nx48830), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48831 (.Y (nx48830), .A0 (ram_255__5), .A1 (nx65606), .S0 (
             nx64354)) ;
    dffr reg_ram_254__5 (.Q (ram_254__5), .QB (\$dummy [1295]), .D (nx48840), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48841 (.Y (nx48840), .A0 (ram_254__5), .A1 (nx65606), .S0 (
             nx64358)) ;
    oai21 ix60059 (.Y (nx60058), .A0 (nx17730), .A1 (nx17652), .B0 (nx65100)) ;
    nand04 ix17731 (.Y (nx17730), .A0 (nx60061), .A1 (nx60069), .A2 (nx60077), .A3 (
           nx60085)) ;
    aoi22 ix60062 (.Y (nx60061), .A0 (ram_224__5), .A1 (nx64510), .B0 (
          ram_225__5), .B1 (nx64548)) ;
    dffr reg_ram_224__5 (.Q (ram_224__5), .QB (\$dummy [1296]), .D (nx48820), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48821 (.Y (nx48820), .A0 (ram_224__5), .A1 (nx65606), .S0 (
             nx64344)) ;
    dffr reg_ram_225__5 (.Q (ram_225__5), .QB (\$dummy [1297]), .D (nx48810), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48811 (.Y (nx48810), .A0 (ram_225__5), .A1 (nx65606), .S0 (
             nx64340)) ;
    aoi22 ix60070 (.Y (nx60069), .A0 (ram_227__5), .A1 (nx64586), .B0 (
          ram_226__5), .B1 (nx64624)) ;
    dffr reg_ram_227__5 (.Q (ram_227__5), .QB (\$dummy [1298]), .D (nx48790), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48791 (.Y (nx48790), .A0 (ram_227__5), .A1 (nx65606), .S0 (
             nx64332)) ;
    dffr reg_ram_226__5 (.Q (ram_226__5), .QB (\$dummy [1299]), .D (nx48800), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48801 (.Y (nx48800), .A0 (ram_226__5), .A1 (nx65606), .S0 (
             nx64336)) ;
    aoi22 ix60078 (.Y (nx60077), .A0 (ram_228__5), .A1 (nx64662), .B0 (
          ram_229__5), .B1 (nx64700)) ;
    dffr reg_ram_228__5 (.Q (ram_228__5), .QB (\$dummy [1300]), .D (nx48780), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48781 (.Y (nx48780), .A0 (ram_228__5), .A1 (nx65606), .S0 (
             nx64328)) ;
    dffr reg_ram_229__5 (.Q (ram_229__5), .QB (\$dummy [1301]), .D (nx48770), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48771 (.Y (nx48770), .A0 (ram_229__5), .A1 (nx65608), .S0 (
             nx64324)) ;
    aoi22 ix60086 (.Y (nx60085), .A0 (ram_231__5), .A1 (nx64738), .B0 (
          ram_230__5), .B1 (nx64776)) ;
    dffr reg_ram_231__5 (.Q (ram_231__5), .QB (\$dummy [1302]), .D (nx48750), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48751 (.Y (nx48750), .A0 (ram_231__5), .A1 (nx65608), .S0 (
             nx64316)) ;
    dffr reg_ram_230__5 (.Q (ram_230__5), .QB (\$dummy [1303]), .D (nx48760), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48761 (.Y (nx48760), .A0 (ram_230__5), .A1 (nx65608), .S0 (
             nx64320)) ;
    nand04 ix17653 (.Y (nx17652), .A0 (nx60094), .A1 (nx60102), .A2 (nx60110), .A3 (
           nx60118)) ;
    aoi22 ix60095 (.Y (nx60094), .A0 (ram_232__5), .A1 (nx64814), .B0 (
          ram_233__5), .B1 (nx64852)) ;
    dffr reg_ram_232__5 (.Q (ram_232__5), .QB (\$dummy [1304]), .D (nx48740), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48741 (.Y (nx48740), .A0 (ram_232__5), .A1 (nx65608), .S0 (
             nx64312)) ;
    dffr reg_ram_233__5 (.Q (ram_233__5), .QB (\$dummy [1305]), .D (nx48730), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48731 (.Y (nx48730), .A0 (ram_233__5), .A1 (nx65608), .S0 (
             nx64308)) ;
    aoi22 ix60103 (.Y (nx60102), .A0 (ram_235__5), .A1 (nx64890), .B0 (
          ram_234__5), .B1 (nx64928)) ;
    dffr reg_ram_235__5 (.Q (ram_235__5), .QB (\$dummy [1306]), .D (nx48710), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48711 (.Y (nx48710), .A0 (ram_235__5), .A1 (nx65608), .S0 (
             nx64300)) ;
    dffr reg_ram_234__5 (.Q (ram_234__5), .QB (\$dummy [1307]), .D (nx48720), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48721 (.Y (nx48720), .A0 (ram_234__5), .A1 (nx65608), .S0 (
             nx64304)) ;
    aoi22 ix60111 (.Y (nx60110), .A0 (ram_236__5), .A1 (nx64966), .B0 (
          ram_237__5), .B1 (nx65004)) ;
    dffr reg_ram_236__5 (.Q (ram_236__5), .QB (\$dummy [1308]), .D (nx48700), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48701 (.Y (nx48700), .A0 (ram_236__5), .A1 (nx65610), .S0 (
             nx64296)) ;
    dffr reg_ram_237__5 (.Q (ram_237__5), .QB (\$dummy [1309]), .D (nx48690), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48691 (.Y (nx48690), .A0 (ram_237__5), .A1 (nx65610), .S0 (
             nx64292)) ;
    aoi22 ix60119 (.Y (nx60118), .A0 (ram_239__5), .A1 (nx65042), .B0 (
          ram_238__5), .B1 (nx65080)) ;
    dffr reg_ram_239__5 (.Q (ram_239__5), .QB (\$dummy [1310]), .D (nx48670), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48671 (.Y (nx48670), .A0 (ram_239__5), .A1 (nx65610), .S0 (
             nx64284)) ;
    dffr reg_ram_238__5 (.Q (ram_238__5), .QB (\$dummy [1311]), .D (nx48680), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48681 (.Y (nx48680), .A0 (ram_238__5), .A1 (nx65610), .S0 (
             nx64288)) ;
    oai21 ix60127 (.Y (nx60126), .A0 (nx17566), .A1 (nx17488), .B0 (nx65104)) ;
    nand04 ix17567 (.Y (nx17566), .A0 (nx60129), .A1 (nx60137), .A2 (nx60145), .A3 (
           nx60153)) ;
    aoi22 ix60130 (.Y (nx60129), .A0 (ram_208__5), .A1 (nx64510), .B0 (
          ram_209__5), .B1 (nx64548)) ;
    dffr reg_ram_208__5 (.Q (ram_208__5), .QB (\$dummy [1312]), .D (nx48660), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48661 (.Y (nx48660), .A0 (ram_208__5), .A1 (nx65610), .S0 (
             nx64274)) ;
    dffr reg_ram_209__5 (.Q (ram_209__5), .QB (\$dummy [1313]), .D (nx48650), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48651 (.Y (nx48650), .A0 (ram_209__5), .A1 (nx65610), .S0 (
             nx64270)) ;
    aoi22 ix60138 (.Y (nx60137), .A0 (ram_211__5), .A1 (nx64586), .B0 (
          ram_210__5), .B1 (nx64624)) ;
    dffr reg_ram_211__5 (.Q (ram_211__5), .QB (\$dummy [1314]), .D (nx48630), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48631 (.Y (nx48630), .A0 (ram_211__5), .A1 (nx65610), .S0 (
             nx64262)) ;
    dffr reg_ram_210__5 (.Q (ram_210__5), .QB (\$dummy [1315]), .D (nx48640), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48641 (.Y (nx48640), .A0 (ram_210__5), .A1 (nx65612), .S0 (
             nx64266)) ;
    aoi22 ix60146 (.Y (nx60145), .A0 (ram_212__5), .A1 (nx64662), .B0 (
          ram_213__5), .B1 (nx64700)) ;
    dffr reg_ram_212__5 (.Q (ram_212__5), .QB (\$dummy [1316]), .D (nx48620), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48621 (.Y (nx48620), .A0 (ram_212__5), .A1 (nx65612), .S0 (
             nx64258)) ;
    dffr reg_ram_213__5 (.Q (ram_213__5), .QB (\$dummy [1317]), .D (nx48610), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48611 (.Y (nx48610), .A0 (ram_213__5), .A1 (nx65612), .S0 (
             nx64254)) ;
    aoi22 ix60154 (.Y (nx60153), .A0 (ram_215__5), .A1 (nx64738), .B0 (
          ram_214__5), .B1 (nx64776)) ;
    dffr reg_ram_215__5 (.Q (ram_215__5), .QB (\$dummy [1318]), .D (nx48590), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48591 (.Y (nx48590), .A0 (ram_215__5), .A1 (nx65612), .S0 (
             nx64246)) ;
    dffr reg_ram_214__5 (.Q (ram_214__5), .QB (\$dummy [1319]), .D (nx48600), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48601 (.Y (nx48600), .A0 (ram_214__5), .A1 (nx65612), .S0 (
             nx64250)) ;
    nand04 ix17489 (.Y (nx17488), .A0 (nx60162), .A1 (nx60170), .A2 (nx60178), .A3 (
           nx60186)) ;
    aoi22 ix60163 (.Y (nx60162), .A0 (ram_216__5), .A1 (nx64814), .B0 (
          ram_217__5), .B1 (nx64852)) ;
    dffr reg_ram_216__5 (.Q (ram_216__5), .QB (\$dummy [1320]), .D (nx48580), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48581 (.Y (nx48580), .A0 (ram_216__5), .A1 (nx65612), .S0 (
             nx64242)) ;
    dffr reg_ram_217__5 (.Q (ram_217__5), .QB (\$dummy [1321]), .D (nx48570), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48571 (.Y (nx48570), .A0 (ram_217__5), .A1 (nx65612), .S0 (
             nx64238)) ;
    aoi22 ix60171 (.Y (nx60170), .A0 (ram_219__5), .A1 (nx64890), .B0 (
          ram_218__5), .B1 (nx64928)) ;
    dffr reg_ram_219__5 (.Q (ram_219__5), .QB (\$dummy [1322]), .D (nx48550), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48551 (.Y (nx48550), .A0 (ram_219__5), .A1 (nx65614), .S0 (
             nx64230)) ;
    dffr reg_ram_218__5 (.Q (ram_218__5), .QB (\$dummy [1323]), .D (nx48560), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48561 (.Y (nx48560), .A0 (ram_218__5), .A1 (nx65614), .S0 (
             nx64234)) ;
    aoi22 ix60179 (.Y (nx60178), .A0 (ram_220__5), .A1 (nx64966), .B0 (
          ram_221__5), .B1 (nx65004)) ;
    dffr reg_ram_220__5 (.Q (ram_220__5), .QB (\$dummy [1324]), .D (nx48540), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48541 (.Y (nx48540), .A0 (ram_220__5), .A1 (nx65614), .S0 (
             nx64226)) ;
    dffr reg_ram_221__5 (.Q (ram_221__5), .QB (\$dummy [1325]), .D (nx48530), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48531 (.Y (nx48530), .A0 (ram_221__5), .A1 (nx65614), .S0 (
             nx64222)) ;
    aoi22 ix60187 (.Y (nx60186), .A0 (ram_223__5), .A1 (nx65042), .B0 (
          ram_222__5), .B1 (nx65080)) ;
    dffr reg_ram_223__5 (.Q (ram_223__5), .QB (\$dummy [1326]), .D (nx48510), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48511 (.Y (nx48510), .A0 (ram_223__5), .A1 (nx65614), .S0 (
             nx64214)) ;
    dffr reg_ram_222__5 (.Q (ram_222__5), .QB (\$dummy [1327]), .D (nx48520), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48521 (.Y (nx48520), .A0 (ram_222__5), .A1 (nx65614), .S0 (
             nx64218)) ;
    oai21 ix60195 (.Y (nx60194), .A0 (nx17404), .A1 (nx17326), .B0 (nx65108)) ;
    nand04 ix17405 (.Y (nx17404), .A0 (nx60197), .A1 (nx60205), .A2 (nx60213), .A3 (
           nx60221)) ;
    aoi22 ix60198 (.Y (nx60197), .A0 (ram_192__5), .A1 (nx64512), .B0 (
          ram_193__5), .B1 (nx64550)) ;
    dffr reg_ram_192__5 (.Q (ram_192__5), .QB (\$dummy [1328]), .D (nx48500), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48501 (.Y (nx48500), .A0 (ram_192__5), .A1 (nx65614), .S0 (
             nx64204)) ;
    dffr reg_ram_193__5 (.Q (ram_193__5), .QB (\$dummy [1329]), .D (nx48490), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48491 (.Y (nx48490), .A0 (ram_193__5), .A1 (nx65616), .S0 (
             nx64200)) ;
    aoi22 ix60206 (.Y (nx60205), .A0 (ram_195__5), .A1 (nx64588), .B0 (
          ram_194__5), .B1 (nx64626)) ;
    dffr reg_ram_195__5 (.Q (ram_195__5), .QB (\$dummy [1330]), .D (nx48470), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48471 (.Y (nx48470), .A0 (ram_195__5), .A1 (nx65616), .S0 (
             nx64192)) ;
    dffr reg_ram_194__5 (.Q (ram_194__5), .QB (\$dummy [1331]), .D (nx48480), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48481 (.Y (nx48480), .A0 (ram_194__5), .A1 (nx65616), .S0 (
             nx64196)) ;
    aoi22 ix60214 (.Y (nx60213), .A0 (ram_196__5), .A1 (nx64664), .B0 (
          ram_197__5), .B1 (nx64702)) ;
    dffr reg_ram_196__5 (.Q (ram_196__5), .QB (\$dummy [1332]), .D (nx48460), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48461 (.Y (nx48460), .A0 (ram_196__5), .A1 (nx65616), .S0 (
             nx64188)) ;
    dffr reg_ram_197__5 (.Q (ram_197__5), .QB (\$dummy [1333]), .D (nx48450), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48451 (.Y (nx48450), .A0 (ram_197__5), .A1 (nx65616), .S0 (
             nx64184)) ;
    aoi22 ix60222 (.Y (nx60221), .A0 (ram_199__5), .A1 (nx64740), .B0 (
          ram_198__5), .B1 (nx64778)) ;
    dffr reg_ram_199__5 (.Q (ram_199__5), .QB (\$dummy [1334]), .D (nx48430), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48431 (.Y (nx48430), .A0 (ram_199__5), .A1 (nx65616), .S0 (
             nx64176)) ;
    dffr reg_ram_198__5 (.Q (ram_198__5), .QB (\$dummy [1335]), .D (nx48440), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48441 (.Y (nx48440), .A0 (ram_198__5), .A1 (nx65616), .S0 (
             nx64180)) ;
    nand04 ix17327 (.Y (nx17326), .A0 (nx60230), .A1 (nx60238), .A2 (nx60246), .A3 (
           nx60254)) ;
    aoi22 ix60231 (.Y (nx60230), .A0 (ram_200__5), .A1 (nx64816), .B0 (
          ram_201__5), .B1 (nx64854)) ;
    dffr reg_ram_200__5 (.Q (ram_200__5), .QB (\$dummy [1336]), .D (nx48420), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48421 (.Y (nx48420), .A0 (ram_200__5), .A1 (nx65618), .S0 (
             nx64172)) ;
    dffr reg_ram_201__5 (.Q (ram_201__5), .QB (\$dummy [1337]), .D (nx48410), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48411 (.Y (nx48410), .A0 (ram_201__5), .A1 (nx65618), .S0 (
             nx64168)) ;
    aoi22 ix60239 (.Y (nx60238), .A0 (ram_203__5), .A1 (nx64892), .B0 (
          ram_202__5), .B1 (nx64930)) ;
    dffr reg_ram_203__5 (.Q (ram_203__5), .QB (\$dummy [1338]), .D (nx48390), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48391 (.Y (nx48390), .A0 (ram_203__5), .A1 (nx65618), .S0 (
             nx64160)) ;
    dffr reg_ram_202__5 (.Q (ram_202__5), .QB (\$dummy [1339]), .D (nx48400), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48401 (.Y (nx48400), .A0 (ram_202__5), .A1 (nx65618), .S0 (
             nx64164)) ;
    aoi22 ix60247 (.Y (nx60246), .A0 (ram_204__5), .A1 (nx64968), .B0 (
          ram_205__5), .B1 (nx65006)) ;
    dffr reg_ram_204__5 (.Q (ram_204__5), .QB (\$dummy [1340]), .D (nx48380), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48381 (.Y (nx48380), .A0 (ram_204__5), .A1 (nx65618), .S0 (
             nx64156)) ;
    dffr reg_ram_205__5 (.Q (ram_205__5), .QB (\$dummy [1341]), .D (nx48370), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48371 (.Y (nx48370), .A0 (ram_205__5), .A1 (nx65618), .S0 (
             nx64152)) ;
    aoi22 ix60255 (.Y (nx60254), .A0 (ram_207__5), .A1 (nx65044), .B0 (
          ram_206__5), .B1 (nx65082)) ;
    dffr reg_ram_207__5 (.Q (ram_207__5), .QB (\$dummy [1342]), .D (nx48350), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48351 (.Y (nx48350), .A0 (ram_207__5), .A1 (nx65618), .S0 (
             nx64144)) ;
    dffr reg_ram_206__5 (.Q (ram_206__5), .QB (\$dummy [1343]), .D (nx48360), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48361 (.Y (nx48360), .A0 (ram_206__5), .A1 (nx65620), .S0 (
             nx64148)) ;
    nand04 ix17249 (.Y (nx17248), .A0 (nx60263), .A1 (nx60331), .A2 (nx60399), .A3 (
           nx60467)) ;
    oai21 ix60264 (.Y (nx60263), .A0 (nx17238), .A1 (nx17160), .B0 (nx65112)) ;
    nand04 ix17239 (.Y (nx17238), .A0 (nx60266), .A1 (nx60274), .A2 (nx60282), .A3 (
           nx60290)) ;
    aoi22 ix60267 (.Y (nx60266), .A0 (ram_80__5), .A1 (nx64512), .B0 (ram_81__5)
          , .B1 (nx64550)) ;
    dffr reg_ram_80__5 (.Q (ram_80__5), .QB (\$dummy [1344]), .D (nx48340), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48341 (.Y (nx48340), .A0 (ram_80__5), .A1 (nx65620), .S0 (nx64134
             )) ;
    dffr reg_ram_81__5 (.Q (ram_81__5), .QB (\$dummy [1345]), .D (nx48330), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48331 (.Y (nx48330), .A0 (ram_81__5), .A1 (nx65620), .S0 (nx64130
             )) ;
    aoi22 ix60275 (.Y (nx60274), .A0 (ram_83__5), .A1 (nx64588), .B0 (ram_82__5)
          , .B1 (nx64626)) ;
    dffr reg_ram_83__5 (.Q (ram_83__5), .QB (\$dummy [1346]), .D (nx48310), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48311 (.Y (nx48310), .A0 (ram_83__5), .A1 (nx65620), .S0 (nx64122
             )) ;
    dffr reg_ram_82__5 (.Q (ram_82__5), .QB (\$dummy [1347]), .D (nx48320), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48321 (.Y (nx48320), .A0 (ram_82__5), .A1 (nx65620), .S0 (nx64126
             )) ;
    aoi22 ix60283 (.Y (nx60282), .A0 (ram_84__5), .A1 (nx64664), .B0 (ram_85__5)
          , .B1 (nx64702)) ;
    dffr reg_ram_84__5 (.Q (ram_84__5), .QB (\$dummy [1348]), .D (nx48300), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48301 (.Y (nx48300), .A0 (ram_84__5), .A1 (nx65620), .S0 (nx64118
             )) ;
    dffr reg_ram_85__5 (.Q (ram_85__5), .QB (\$dummy [1349]), .D (nx48290), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48291 (.Y (nx48290), .A0 (ram_85__5), .A1 (nx65620), .S0 (nx64114
             )) ;
    aoi22 ix60291 (.Y (nx60290), .A0 (ram_87__5), .A1 (nx64740), .B0 (ram_86__5)
          , .B1 (nx64778)) ;
    dffr reg_ram_87__5 (.Q (ram_87__5), .QB (\$dummy [1350]), .D (nx48270), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48271 (.Y (nx48270), .A0 (ram_87__5), .A1 (nx65622), .S0 (nx64106
             )) ;
    dffr reg_ram_86__5 (.Q (ram_86__5), .QB (\$dummy [1351]), .D (nx48280), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48281 (.Y (nx48280), .A0 (ram_86__5), .A1 (nx65622), .S0 (nx64110
             )) ;
    nand04 ix17161 (.Y (nx17160), .A0 (nx60299), .A1 (nx60307), .A2 (nx60315), .A3 (
           nx60323)) ;
    aoi22 ix60300 (.Y (nx60299), .A0 (ram_88__5), .A1 (nx64816), .B0 (ram_89__5)
          , .B1 (nx64854)) ;
    dffr reg_ram_88__5 (.Q (ram_88__5), .QB (\$dummy [1352]), .D (nx48260), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48261 (.Y (nx48260), .A0 (ram_88__5), .A1 (nx65622), .S0 (nx64102
             )) ;
    dffr reg_ram_89__5 (.Q (ram_89__5), .QB (\$dummy [1353]), .D (nx48250), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48251 (.Y (nx48250), .A0 (ram_89__5), .A1 (nx65622), .S0 (nx64098
             )) ;
    aoi22 ix60308 (.Y (nx60307), .A0 (ram_91__5), .A1 (nx64892), .B0 (ram_90__5)
          , .B1 (nx64930)) ;
    dffr reg_ram_91__5 (.Q (ram_91__5), .QB (\$dummy [1354]), .D (nx48230), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48231 (.Y (nx48230), .A0 (ram_91__5), .A1 (nx65622), .S0 (nx64090
             )) ;
    dffr reg_ram_90__5 (.Q (ram_90__5), .QB (\$dummy [1355]), .D (nx48240), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48241 (.Y (nx48240), .A0 (ram_90__5), .A1 (nx65622), .S0 (nx64094
             )) ;
    aoi22 ix60316 (.Y (nx60315), .A0 (ram_92__5), .A1 (nx64968), .B0 (ram_93__5)
          , .B1 (nx65006)) ;
    dffr reg_ram_92__5 (.Q (ram_92__5), .QB (\$dummy [1356]), .D (nx48220), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48221 (.Y (nx48220), .A0 (ram_92__5), .A1 (nx65622), .S0 (nx64086
             )) ;
    dffr reg_ram_93__5 (.Q (ram_93__5), .QB (\$dummy [1357]), .D (nx48210), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48211 (.Y (nx48210), .A0 (ram_93__5), .A1 (nx65624), .S0 (nx64082
             )) ;
    aoi22 ix60324 (.Y (nx60323), .A0 (ram_95__5), .A1 (nx65044), .B0 (ram_94__5)
          , .B1 (nx65082)) ;
    dffr reg_ram_95__5 (.Q (ram_95__5), .QB (\$dummy [1358]), .D (nx48190), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48191 (.Y (nx48190), .A0 (ram_95__5), .A1 (nx65624), .S0 (nx64074
             )) ;
    dffr reg_ram_94__5 (.Q (ram_94__5), .QB (\$dummy [1359]), .D (nx48200), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48201 (.Y (nx48200), .A0 (ram_94__5), .A1 (nx65624), .S0 (nx64078
             )) ;
    oai21 ix60332 (.Y (nx60331), .A0 (nx17076), .A1 (nx16998), .B0 (nx65116)) ;
    nand04 ix17077 (.Y (nx17076), .A0 (nx60334), .A1 (nx60342), .A2 (nx60350), .A3 (
           nx60358)) ;
    aoi22 ix60335 (.Y (nx60334), .A0 (ram_64__5), .A1 (nx64512), .B0 (ram_65__5)
          , .B1 (nx64550)) ;
    dffr reg_ram_64__5 (.Q (ram_64__5), .QB (\$dummy [1360]), .D (nx48180), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48181 (.Y (nx48180), .A0 (ram_64__5), .A1 (nx65624), .S0 (nx64064
             )) ;
    dffr reg_ram_65__5 (.Q (ram_65__5), .QB (\$dummy [1361]), .D (nx48170), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48171 (.Y (nx48170), .A0 (ram_65__5), .A1 (nx65624), .S0 (nx64060
             )) ;
    aoi22 ix60343 (.Y (nx60342), .A0 (ram_67__5), .A1 (nx64588), .B0 (ram_66__5)
          , .B1 (nx64626)) ;
    dffr reg_ram_67__5 (.Q (ram_67__5), .QB (\$dummy [1362]), .D (nx48150), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48151 (.Y (nx48150), .A0 (ram_67__5), .A1 (nx65624), .S0 (nx64052
             )) ;
    dffr reg_ram_66__5 (.Q (ram_66__5), .QB (\$dummy [1363]), .D (nx48160), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48161 (.Y (nx48160), .A0 (ram_66__5), .A1 (nx65624), .S0 (nx64056
             )) ;
    aoi22 ix60351 (.Y (nx60350), .A0 (ram_68__5), .A1 (nx64664), .B0 (ram_69__5)
          , .B1 (nx64702)) ;
    dffr reg_ram_68__5 (.Q (ram_68__5), .QB (\$dummy [1364]), .D (nx48140), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48141 (.Y (nx48140), .A0 (ram_68__5), .A1 (nx65626), .S0 (nx64048
             )) ;
    dffr reg_ram_69__5 (.Q (ram_69__5), .QB (\$dummy [1365]), .D (nx48130), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48131 (.Y (nx48130), .A0 (ram_69__5), .A1 (nx65626), .S0 (nx64044
             )) ;
    aoi22 ix60359 (.Y (nx60358), .A0 (ram_71__5), .A1 (nx64740), .B0 (ram_70__5)
          , .B1 (nx64778)) ;
    dffr reg_ram_71__5 (.Q (ram_71__5), .QB (\$dummy [1366]), .D (nx48110), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48111 (.Y (nx48110), .A0 (ram_71__5), .A1 (nx65626), .S0 (nx64036
             )) ;
    dffr reg_ram_70__5 (.Q (ram_70__5), .QB (\$dummy [1367]), .D (nx48120), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48121 (.Y (nx48120), .A0 (ram_70__5), .A1 (nx65626), .S0 (nx64040
             )) ;
    nand04 ix16999 (.Y (nx16998), .A0 (nx60367), .A1 (nx60375), .A2 (nx60383), .A3 (
           nx60391)) ;
    aoi22 ix60368 (.Y (nx60367), .A0 (ram_72__5), .A1 (nx64816), .B0 (ram_73__5)
          , .B1 (nx64854)) ;
    dffr reg_ram_72__5 (.Q (ram_72__5), .QB (\$dummy [1368]), .D (nx48100), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48101 (.Y (nx48100), .A0 (ram_72__5), .A1 (nx65626), .S0 (nx64032
             )) ;
    dffr reg_ram_73__5 (.Q (ram_73__5), .QB (\$dummy [1369]), .D (nx48090), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48091 (.Y (nx48090), .A0 (ram_73__5), .A1 (nx65626), .S0 (nx64028
             )) ;
    aoi22 ix60376 (.Y (nx60375), .A0 (ram_75__5), .A1 (nx64892), .B0 (ram_74__5)
          , .B1 (nx64930)) ;
    dffr reg_ram_75__5 (.Q (ram_75__5), .QB (\$dummy [1370]), .D (nx48070), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48071 (.Y (nx48070), .A0 (ram_75__5), .A1 (nx65626), .S0 (nx64020
             )) ;
    dffr reg_ram_74__5 (.Q (ram_74__5), .QB (\$dummy [1371]), .D (nx48080), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48081 (.Y (nx48080), .A0 (ram_74__5), .A1 (nx65628), .S0 (nx64024
             )) ;
    aoi22 ix60384 (.Y (nx60383), .A0 (ram_76__5), .A1 (nx64968), .B0 (ram_77__5)
          , .B1 (nx65006)) ;
    dffr reg_ram_76__5 (.Q (ram_76__5), .QB (\$dummy [1372]), .D (nx48060), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48061 (.Y (nx48060), .A0 (ram_76__5), .A1 (nx65628), .S0 (nx64016
             )) ;
    dffr reg_ram_77__5 (.Q (ram_77__5), .QB (\$dummy [1373]), .D (nx48050), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48051 (.Y (nx48050), .A0 (ram_77__5), .A1 (nx65628), .S0 (nx64012
             )) ;
    aoi22 ix60392 (.Y (nx60391), .A0 (ram_79__5), .A1 (nx65044), .B0 (ram_78__5)
          , .B1 (nx65082)) ;
    dffr reg_ram_79__5 (.Q (ram_79__5), .QB (\$dummy [1374]), .D (nx48030), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48031 (.Y (nx48030), .A0 (ram_79__5), .A1 (nx65628), .S0 (nx64004
             )) ;
    dffr reg_ram_78__5 (.Q (ram_78__5), .QB (\$dummy [1375]), .D (nx48040), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48041 (.Y (nx48040), .A0 (ram_78__5), .A1 (nx65628), .S0 (nx64008
             )) ;
    oai21 ix60400 (.Y (nx60399), .A0 (nx16912), .A1 (nx16834), .B0 (nx65120)) ;
    nand04 ix16913 (.Y (nx16912), .A0 (nx60402), .A1 (nx60410), .A2 (nx60418), .A3 (
           nx60426)) ;
    aoi22 ix60403 (.Y (nx60402), .A0 (ram_48__5), .A1 (nx64512), .B0 (ram_49__5)
          , .B1 (nx64550)) ;
    dffr reg_ram_48__5 (.Q (ram_48__5), .QB (\$dummy [1376]), .D (nx48020), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48021 (.Y (nx48020), .A0 (ram_48__5), .A1 (nx65628), .S0 (nx63994
             )) ;
    dffr reg_ram_49__5 (.Q (ram_49__5), .QB (\$dummy [1377]), .D (nx48010), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48011 (.Y (nx48010), .A0 (ram_49__5), .A1 (nx65628), .S0 (nx63990
             )) ;
    aoi22 ix60411 (.Y (nx60410), .A0 (ram_51__5), .A1 (nx64588), .B0 (ram_50__5)
          , .B1 (nx64626)) ;
    dffr reg_ram_51__5 (.Q (ram_51__5), .QB (\$dummy [1378]), .D (nx47990), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47991 (.Y (nx47990), .A0 (ram_51__5), .A1 (nx65630), .S0 (nx63982
             )) ;
    dffr reg_ram_50__5 (.Q (ram_50__5), .QB (\$dummy [1379]), .D (nx48000), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48001 (.Y (nx48000), .A0 (ram_50__5), .A1 (nx65630), .S0 (nx63986
             )) ;
    aoi22 ix60419 (.Y (nx60418), .A0 (ram_52__5), .A1 (nx64664), .B0 (ram_53__5)
          , .B1 (nx64702)) ;
    dffr reg_ram_52__5 (.Q (ram_52__5), .QB (\$dummy [1380]), .D (nx47980), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47981 (.Y (nx47980), .A0 (ram_52__5), .A1 (nx65630), .S0 (nx63978
             )) ;
    dffr reg_ram_53__5 (.Q (ram_53__5), .QB (\$dummy [1381]), .D (nx47970), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47971 (.Y (nx47970), .A0 (ram_53__5), .A1 (nx65630), .S0 (nx63974
             )) ;
    aoi22 ix60427 (.Y (nx60426), .A0 (ram_55__5), .A1 (nx64740), .B0 (ram_54__5)
          , .B1 (nx64778)) ;
    dffr reg_ram_55__5 (.Q (ram_55__5), .QB (\$dummy [1382]), .D (nx47950), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47951 (.Y (nx47950), .A0 (ram_55__5), .A1 (nx65630), .S0 (nx63966
             )) ;
    dffr reg_ram_54__5 (.Q (ram_54__5), .QB (\$dummy [1383]), .D (nx47960), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47961 (.Y (nx47960), .A0 (ram_54__5), .A1 (nx65630), .S0 (nx63970
             )) ;
    nand04 ix16835 (.Y (nx16834), .A0 (nx60435), .A1 (nx60443), .A2 (nx60451), .A3 (
           nx60459)) ;
    aoi22 ix60436 (.Y (nx60435), .A0 (ram_56__5), .A1 (nx64816), .B0 (ram_57__5)
          , .B1 (nx64854)) ;
    dffr reg_ram_56__5 (.Q (ram_56__5), .QB (\$dummy [1384]), .D (nx47940), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47941 (.Y (nx47940), .A0 (ram_56__5), .A1 (nx65630), .S0 (nx63962
             )) ;
    dffr reg_ram_57__5 (.Q (ram_57__5), .QB (\$dummy [1385]), .D (nx47930), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47931 (.Y (nx47930), .A0 (ram_57__5), .A1 (nx65632), .S0 (nx63958
             )) ;
    aoi22 ix60444 (.Y (nx60443), .A0 (ram_59__5), .A1 (nx64892), .B0 (ram_58__5)
          , .B1 (nx64930)) ;
    dffr reg_ram_59__5 (.Q (ram_59__5), .QB (\$dummy [1386]), .D (nx47910), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47911 (.Y (nx47910), .A0 (ram_59__5), .A1 (nx65632), .S0 (nx63950
             )) ;
    dffr reg_ram_58__5 (.Q (ram_58__5), .QB (\$dummy [1387]), .D (nx47920), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47921 (.Y (nx47920), .A0 (ram_58__5), .A1 (nx65632), .S0 (nx63954
             )) ;
    aoi22 ix60452 (.Y (nx60451), .A0 (ram_60__5), .A1 (nx64968), .B0 (ram_61__5)
          , .B1 (nx65006)) ;
    dffr reg_ram_60__5 (.Q (ram_60__5), .QB (\$dummy [1388]), .D (nx47900), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47901 (.Y (nx47900), .A0 (ram_60__5), .A1 (nx65632), .S0 (nx63946
             )) ;
    dffr reg_ram_61__5 (.Q (ram_61__5), .QB (\$dummy [1389]), .D (nx47890), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47891 (.Y (nx47890), .A0 (ram_61__5), .A1 (nx65632), .S0 (nx63942
             )) ;
    aoi22 ix60460 (.Y (nx60459), .A0 (ram_63__5), .A1 (nx65044), .B0 (ram_62__5)
          , .B1 (nx65082)) ;
    dffr reg_ram_63__5 (.Q (ram_63__5), .QB (\$dummy [1390]), .D (nx47870), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47871 (.Y (nx47870), .A0 (ram_63__5), .A1 (nx65632), .S0 (nx63934
             )) ;
    dffr reg_ram_62__5 (.Q (ram_62__5), .QB (\$dummy [1391]), .D (nx47880), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47881 (.Y (nx47880), .A0 (ram_62__5), .A1 (nx65632), .S0 (nx63938
             )) ;
    oai21 ix60468 (.Y (nx60467), .A0 (nx16750), .A1 (nx16672), .B0 (nx65124)) ;
    nand04 ix16751 (.Y (nx16750), .A0 (nx60470), .A1 (nx60478), .A2 (nx60486), .A3 (
           nx60494)) ;
    aoi22 ix60471 (.Y (nx60470), .A0 (ram_32__5), .A1 (nx64512), .B0 (ram_33__5)
          , .B1 (nx64550)) ;
    dffr reg_ram_32__5 (.Q (ram_32__5), .QB (\$dummy [1392]), .D (nx47860), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47861 (.Y (nx47860), .A0 (ram_32__5), .A1 (nx65634), .S0 (nx63924
             )) ;
    dffr reg_ram_33__5 (.Q (ram_33__5), .QB (\$dummy [1393]), .D (nx47850), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47851 (.Y (nx47850), .A0 (ram_33__5), .A1 (nx65634), .S0 (nx63920
             )) ;
    aoi22 ix60479 (.Y (nx60478), .A0 (ram_35__5), .A1 (nx64588), .B0 (ram_34__5)
          , .B1 (nx64626)) ;
    dffr reg_ram_35__5 (.Q (ram_35__5), .QB (\$dummy [1394]), .D (nx47830), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47831 (.Y (nx47830), .A0 (ram_35__5), .A1 (nx65634), .S0 (nx63912
             )) ;
    dffr reg_ram_34__5 (.Q (ram_34__5), .QB (\$dummy [1395]), .D (nx47840), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47841 (.Y (nx47840), .A0 (ram_34__5), .A1 (nx65634), .S0 (nx63916
             )) ;
    aoi22 ix60487 (.Y (nx60486), .A0 (ram_36__5), .A1 (nx64664), .B0 (ram_37__5)
          , .B1 (nx64702)) ;
    dffr reg_ram_36__5 (.Q (ram_36__5), .QB (\$dummy [1396]), .D (nx47820), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47821 (.Y (nx47820), .A0 (ram_36__5), .A1 (nx65634), .S0 (nx63908
             )) ;
    dffr reg_ram_37__5 (.Q (ram_37__5), .QB (\$dummy [1397]), .D (nx47810), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47811 (.Y (nx47810), .A0 (ram_37__5), .A1 (nx65634), .S0 (nx63904
             )) ;
    aoi22 ix60495 (.Y (nx60494), .A0 (ram_39__5), .A1 (nx64740), .B0 (ram_38__5)
          , .B1 (nx64778)) ;
    dffr reg_ram_39__5 (.Q (ram_39__5), .QB (\$dummy [1398]), .D (nx47790), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47791 (.Y (nx47790), .A0 (ram_39__5), .A1 (nx65634), .S0 (nx63896
             )) ;
    dffr reg_ram_38__5 (.Q (ram_38__5), .QB (\$dummy [1399]), .D (nx47800), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47801 (.Y (nx47800), .A0 (ram_38__5), .A1 (nx65636), .S0 (nx63900
             )) ;
    nand04 ix16673 (.Y (nx16672), .A0 (nx60503), .A1 (nx60511), .A2 (nx60519), .A3 (
           nx60527)) ;
    aoi22 ix60504 (.Y (nx60503), .A0 (ram_40__5), .A1 (nx64816), .B0 (ram_41__5)
          , .B1 (nx64854)) ;
    dffr reg_ram_40__5 (.Q (ram_40__5), .QB (\$dummy [1400]), .D (nx47780), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47781 (.Y (nx47780), .A0 (ram_40__5), .A1 (nx65636), .S0 (nx63892
             )) ;
    dffr reg_ram_41__5 (.Q (ram_41__5), .QB (\$dummy [1401]), .D (nx47770), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47771 (.Y (nx47770), .A0 (ram_41__5), .A1 (nx65636), .S0 (nx63888
             )) ;
    aoi22 ix60512 (.Y (nx60511), .A0 (ram_43__5), .A1 (nx64892), .B0 (ram_42__5)
          , .B1 (nx64930)) ;
    dffr reg_ram_43__5 (.Q (ram_43__5), .QB (\$dummy [1402]), .D (nx47750), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47751 (.Y (nx47750), .A0 (ram_43__5), .A1 (nx65636), .S0 (nx63880
             )) ;
    dffr reg_ram_42__5 (.Q (ram_42__5), .QB (\$dummy [1403]), .D (nx47760), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47761 (.Y (nx47760), .A0 (ram_42__5), .A1 (nx65636), .S0 (nx63884
             )) ;
    aoi22 ix60520 (.Y (nx60519), .A0 (ram_44__5), .A1 (nx64968), .B0 (ram_45__5)
          , .B1 (nx65006)) ;
    dffr reg_ram_44__5 (.Q (ram_44__5), .QB (\$dummy [1404]), .D (nx47740), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47741 (.Y (nx47740), .A0 (ram_44__5), .A1 (nx65636), .S0 (nx63876
             )) ;
    dffr reg_ram_45__5 (.Q (ram_45__5), .QB (\$dummy [1405]), .D (nx47730), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47731 (.Y (nx47730), .A0 (ram_45__5), .A1 (nx65636), .S0 (nx63872
             )) ;
    aoi22 ix60528 (.Y (nx60527), .A0 (ram_47__5), .A1 (nx65044), .B0 (ram_46__5)
          , .B1 (nx65082)) ;
    dffr reg_ram_47__5 (.Q (ram_47__5), .QB (\$dummy [1406]), .D (nx47710), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47711 (.Y (nx47710), .A0 (ram_47__5), .A1 (nx65638), .S0 (nx63864
             )) ;
    dffr reg_ram_46__5 (.Q (ram_46__5), .QB (\$dummy [1407]), .D (nx47720), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47721 (.Y (nx47720), .A0 (ram_46__5), .A1 (nx65638), .S0 (nx63868
             )) ;
    nand04 ix16593 (.Y (nx16592), .A0 (nx60536), .A1 (nx60604), .A2 (nx60672), .A3 (
           nx60740)) ;
    oai21 ix60537 (.Y (nx60536), .A0 (nx16582), .A1 (nx16504), .B0 (nx65128)) ;
    nand04 ix16583 (.Y (nx16582), .A0 (nx60539), .A1 (nx60547), .A2 (nx60555), .A3 (
           nx60563)) ;
    aoi22 ix60540 (.Y (nx60539), .A0 (ram_16__5), .A1 (nx64512), .B0 (ram_17__5)
          , .B1 (nx64550)) ;
    dffr reg_ram_16__5 (.Q (ram_16__5), .QB (\$dummy [1408]), .D (nx47700), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47701 (.Y (nx47700), .A0 (ram_16__5), .A1 (nx65638), .S0 (nx63854
             )) ;
    dffr reg_ram_17__5 (.Q (ram_17__5), .QB (\$dummy [1409]), .D (nx47690), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47691 (.Y (nx47690), .A0 (ram_17__5), .A1 (nx65638), .S0 (nx63850
             )) ;
    aoi22 ix60548 (.Y (nx60547), .A0 (ram_19__5), .A1 (nx64588), .B0 (ram_18__5)
          , .B1 (nx64626)) ;
    dffr reg_ram_19__5 (.Q (ram_19__5), .QB (\$dummy [1410]), .D (nx47670), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47671 (.Y (nx47670), .A0 (ram_19__5), .A1 (nx65638), .S0 (nx63842
             )) ;
    dffr reg_ram_18__5 (.Q (ram_18__5), .QB (\$dummy [1411]), .D (nx47680), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47681 (.Y (nx47680), .A0 (ram_18__5), .A1 (nx65638), .S0 (nx63846
             )) ;
    aoi22 ix60556 (.Y (nx60555), .A0 (ram_20__5), .A1 (nx64664), .B0 (ram_21__5)
          , .B1 (nx64702)) ;
    dffr reg_ram_20__5 (.Q (ram_20__5), .QB (\$dummy [1412]), .D (nx47660), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47661 (.Y (nx47660), .A0 (ram_20__5), .A1 (nx65638), .S0 (nx63838
             )) ;
    dffr reg_ram_21__5 (.Q (ram_21__5), .QB (\$dummy [1413]), .D (nx47650), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47651 (.Y (nx47650), .A0 (ram_21__5), .A1 (nx65640), .S0 (nx63834
             )) ;
    aoi22 ix60564 (.Y (nx60563), .A0 (ram_23__5), .A1 (nx64740), .B0 (ram_22__5)
          , .B1 (nx64778)) ;
    dffr reg_ram_23__5 (.Q (ram_23__5), .QB (\$dummy [1414]), .D (nx47630), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47631 (.Y (nx47630), .A0 (ram_23__5), .A1 (nx65640), .S0 (nx63826
             )) ;
    dffr reg_ram_22__5 (.Q (ram_22__5), .QB (\$dummy [1415]), .D (nx47640), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47641 (.Y (nx47640), .A0 (ram_22__5), .A1 (nx65640), .S0 (nx63830
             )) ;
    nand04 ix16505 (.Y (nx16504), .A0 (nx60572), .A1 (nx60580), .A2 (nx60588), .A3 (
           nx60596)) ;
    aoi22 ix60573 (.Y (nx60572), .A0 (ram_24__5), .A1 (nx64816), .B0 (ram_25__5)
          , .B1 (nx64854)) ;
    dffr reg_ram_24__5 (.Q (ram_24__5), .QB (\$dummy [1416]), .D (nx47620), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47621 (.Y (nx47620), .A0 (ram_24__5), .A1 (nx65640), .S0 (nx63822
             )) ;
    dffr reg_ram_25__5 (.Q (ram_25__5), .QB (\$dummy [1417]), .D (nx47610), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47611 (.Y (nx47610), .A0 (ram_25__5), .A1 (nx65640), .S0 (nx63818
             )) ;
    aoi22 ix60581 (.Y (nx60580), .A0 (ram_27__5), .A1 (nx64892), .B0 (ram_26__5)
          , .B1 (nx64930)) ;
    dffr reg_ram_27__5 (.Q (ram_27__5), .QB (\$dummy [1418]), .D (nx47590), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47591 (.Y (nx47590), .A0 (ram_27__5), .A1 (nx65640), .S0 (nx63810
             )) ;
    dffr reg_ram_26__5 (.Q (ram_26__5), .QB (\$dummy [1419]), .D (nx47600), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47601 (.Y (nx47600), .A0 (ram_26__5), .A1 (nx65640), .S0 (nx63814
             )) ;
    aoi22 ix60589 (.Y (nx60588), .A0 (ram_28__5), .A1 (nx64968), .B0 (ram_29__5)
          , .B1 (nx65006)) ;
    dffr reg_ram_28__5 (.Q (ram_28__5), .QB (\$dummy [1420]), .D (nx47580), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47581 (.Y (nx47580), .A0 (ram_28__5), .A1 (nx65642), .S0 (nx63806
             )) ;
    dffr reg_ram_29__5 (.Q (ram_29__5), .QB (\$dummy [1421]), .D (nx47570), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47571 (.Y (nx47570), .A0 (ram_29__5), .A1 (nx65642), .S0 (nx63802
             )) ;
    aoi22 ix60597 (.Y (nx60596), .A0 (ram_31__5), .A1 (nx65044), .B0 (ram_30__5)
          , .B1 (nx65082)) ;
    dffr reg_ram_31__5 (.Q (ram_31__5), .QB (\$dummy [1422]), .D (nx47550), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47551 (.Y (nx47550), .A0 (ram_31__5), .A1 (nx65642), .S0 (nx63794
             )) ;
    dffr reg_ram_30__5 (.Q (ram_30__5), .QB (\$dummy [1423]), .D (nx47560), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47561 (.Y (nx47560), .A0 (ram_30__5), .A1 (nx65642), .S0 (nx63798
             )) ;
    oai21 ix60605 (.Y (nx60604), .A0 (nx16420), .A1 (nx16342), .B0 (nx65144)) ;
    nand04 ix16421 (.Y (nx16420), .A0 (nx60607), .A1 (nx60615), .A2 (nx60623), .A3 (
           nx60631)) ;
    aoi22 ix60608 (.Y (nx60607), .A0 (ram_0__5), .A1 (nx64512), .B0 (ram_1__5), 
          .B1 (nx64550)) ;
    dffr reg_ram_0__5 (.Q (ram_0__5), .QB (\$dummy [1424]), .D (nx47540), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47541 (.Y (nx47540), .A0 (nx65642), .A1 (ram_0__5), .S0 (nx65132)
             ) ;
    dffr reg_ram_1__5 (.Q (ram_1__5), .QB (\$dummy [1425]), .D (nx47530), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47531 (.Y (nx47530), .A0 (nx65642), .A1 (ram_1__5), .S0 (nx65146)
             ) ;
    aoi22 ix60616 (.Y (nx60615), .A0 (ram_3__5), .A1 (nx64588), .B0 (ram_2__5), 
          .B1 (nx64626)) ;
    dffr reg_ram_3__5 (.Q (ram_3__5), .QB (\$dummy [1426]), .D (nx47510), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47511 (.Y (nx47510), .A0 (nx65642), .A1 (ram_3__5), .S0 (nx65150)
             ) ;
    dffr reg_ram_2__5 (.Q (ram_2__5), .QB (\$dummy [1427]), .D (nx47520), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47521 (.Y (nx47520), .A0 (nx65644), .A1 (ram_2__5), .S0 (nx65154)
             ) ;
    aoi22 ix60624 (.Y (nx60623), .A0 (ram_4__5), .A1 (nx64664), .B0 (ram_5__5), 
          .B1 (nx64702)) ;
    dffr reg_ram_4__5 (.Q (ram_4__5), .QB (\$dummy [1428]), .D (nx47500), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47501 (.Y (nx47500), .A0 (nx65644), .A1 (ram_4__5), .S0 (nx65158)
             ) ;
    dffr reg_ram_5__5 (.Q (ram_5__5), .QB (\$dummy [1429]), .D (nx47490), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47491 (.Y (nx47490), .A0 (nx65644), .A1 (ram_5__5), .S0 (nx65162)
             ) ;
    aoi22 ix60632 (.Y (nx60631), .A0 (ram_7__5), .A1 (nx64740), .B0 (ram_6__5), 
          .B1 (nx64778)) ;
    dffr reg_ram_7__5 (.Q (ram_7__5), .QB (\$dummy [1430]), .D (nx47470), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47471 (.Y (nx47470), .A0 (nx65644), .A1 (ram_7__5), .S0 (nx65166)
             ) ;
    dffr reg_ram_6__5 (.Q (ram_6__5), .QB (\$dummy [1431]), .D (nx47480), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47481 (.Y (nx47480), .A0 (nx65644), .A1 (ram_6__5), .S0 (nx65170)
             ) ;
    nand04 ix16343 (.Y (nx16342), .A0 (nx60640), .A1 (nx60648), .A2 (nx60656), .A3 (
           nx60664)) ;
    aoi22 ix60641 (.Y (nx60640), .A0 (ram_8__5), .A1 (nx64816), .B0 (ram_9__5), 
          .B1 (nx64854)) ;
    dffr reg_ram_8__5 (.Q (ram_8__5), .QB (\$dummy [1432]), .D (nx47460), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47461 (.Y (nx47460), .A0 (nx65644), .A1 (ram_8__5), .S0 (nx65174)
             ) ;
    dffr reg_ram_9__5 (.Q (ram_9__5), .QB (\$dummy [1433]), .D (nx47450), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47451 (.Y (nx47450), .A0 (nx65644), .A1 (ram_9__5), .S0 (nx65178)
             ) ;
    aoi22 ix60649 (.Y (nx60648), .A0 (ram_11__5), .A1 (nx64892), .B0 (ram_10__5)
          , .B1 (nx64930)) ;
    dffr reg_ram_11__5 (.Q (ram_11__5), .QB (\$dummy [1434]), .D (nx47430), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47431 (.Y (nx47430), .A0 (nx65646), .A1 (ram_11__5), .S0 (nx65182
             )) ;
    dffr reg_ram_10__5 (.Q (ram_10__5), .QB (\$dummy [1435]), .D (nx47440), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47441 (.Y (nx47440), .A0 (nx65646), .A1 (ram_10__5), .S0 (nx65186
             )) ;
    aoi22 ix60657 (.Y (nx60656), .A0 (ram_12__5), .A1 (nx64968), .B0 (ram_13__5)
          , .B1 (nx65006)) ;
    dffr reg_ram_12__5 (.Q (ram_12__5), .QB (\$dummy [1436]), .D (nx47420), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47421 (.Y (nx47420), .A0 (nx65646), .A1 (ram_12__5), .S0 (nx65190
             )) ;
    dffr reg_ram_13__5 (.Q (ram_13__5), .QB (\$dummy [1437]), .D (nx47410), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47411 (.Y (nx47410), .A0 (nx65646), .A1 (ram_13__5), .S0 (nx65194
             )) ;
    aoi22 ix60665 (.Y (nx60664), .A0 (ram_15__5), .A1 (nx65044), .B0 (ram_14__5)
          , .B1 (nx65082)) ;
    dffr reg_ram_15__5 (.Q (ram_15__5), .QB (\$dummy [1438]), .D (nx47390), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47391 (.Y (nx47390), .A0 (nx65646), .A1 (ram_15__5), .S0 (nx65198
             )) ;
    dffr reg_ram_14__5 (.Q (ram_14__5), .QB (\$dummy [1439]), .D (nx47400), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47401 (.Y (nx47400), .A0 (nx65646), .A1 (ram_14__5), .S0 (nx65202
             )) ;
    oai21 ix60673 (.Y (nx60672), .A0 (nx16256), .A1 (nx16178), .B0 (nx65206)) ;
    nand04 ix16257 (.Y (nx16256), .A0 (nx60675), .A1 (nx60683), .A2 (nx60691), .A3 (
           nx60699)) ;
    aoi22 ix60676 (.Y (nx60675), .A0 (ram_96__5), .A1 (nx64514), .B0 (ram_97__5)
          , .B1 (nx64552)) ;
    dffr reg_ram_96__5 (.Q (ram_96__5), .QB (\$dummy [1440]), .D (nx47380), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47381 (.Y (nx47380), .A0 (ram_96__5), .A1 (nx65646), .S0 (nx63784
             )) ;
    dffr reg_ram_97__5 (.Q (ram_97__5), .QB (\$dummy [1441]), .D (nx47370), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47371 (.Y (nx47370), .A0 (ram_97__5), .A1 (nx65648), .S0 (nx63780
             )) ;
    aoi22 ix60684 (.Y (nx60683), .A0 (ram_99__5), .A1 (nx64590), .B0 (ram_98__5)
          , .B1 (nx64628)) ;
    dffr reg_ram_99__5 (.Q (ram_99__5), .QB (\$dummy [1442]), .D (nx47350), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47351 (.Y (nx47350), .A0 (ram_99__5), .A1 (nx65648), .S0 (nx63772
             )) ;
    dffr reg_ram_98__5 (.Q (ram_98__5), .QB (\$dummy [1443]), .D (nx47360), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47361 (.Y (nx47360), .A0 (ram_98__5), .A1 (nx65648), .S0 (nx63776
             )) ;
    aoi22 ix60692 (.Y (nx60691), .A0 (ram_100__5), .A1 (nx64666), .B0 (
          ram_101__5), .B1 (nx64704)) ;
    dffr reg_ram_100__5 (.Q (ram_100__5), .QB (\$dummy [1444]), .D (nx47340), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47341 (.Y (nx47340), .A0 (ram_100__5), .A1 (nx65648), .S0 (
             nx63768)) ;
    dffr reg_ram_101__5 (.Q (ram_101__5), .QB (\$dummy [1445]), .D (nx47330), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47331 (.Y (nx47330), .A0 (ram_101__5), .A1 (nx65648), .S0 (
             nx63764)) ;
    aoi22 ix60700 (.Y (nx60699), .A0 (ram_103__5), .A1 (nx64742), .B0 (
          ram_102__5), .B1 (nx64780)) ;
    dffr reg_ram_103__5 (.Q (ram_103__5), .QB (\$dummy [1446]), .D (nx47310), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47311 (.Y (nx47310), .A0 (ram_103__5), .A1 (nx65648), .S0 (
             nx63756)) ;
    dffr reg_ram_102__5 (.Q (ram_102__5), .QB (\$dummy [1447]), .D (nx47320), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47321 (.Y (nx47320), .A0 (ram_102__5), .A1 (nx65648), .S0 (
             nx63760)) ;
    nand04 ix16179 (.Y (nx16178), .A0 (nx60708), .A1 (nx60716), .A2 (nx60724), .A3 (
           nx60732)) ;
    aoi22 ix60709 (.Y (nx60708), .A0 (ram_104__5), .A1 (nx64818), .B0 (
          ram_105__5), .B1 (nx64856)) ;
    dffr reg_ram_104__5 (.Q (ram_104__5), .QB (\$dummy [1448]), .D (nx47300), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47301 (.Y (nx47300), .A0 (ram_104__5), .A1 (nx65650), .S0 (
             nx63752)) ;
    dffr reg_ram_105__5 (.Q (ram_105__5), .QB (\$dummy [1449]), .D (nx47290), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47291 (.Y (nx47290), .A0 (ram_105__5), .A1 (nx65650), .S0 (
             nx63748)) ;
    aoi22 ix60717 (.Y (nx60716), .A0 (ram_107__5), .A1 (nx64894), .B0 (
          ram_106__5), .B1 (nx64932)) ;
    dffr reg_ram_107__5 (.Q (ram_107__5), .QB (\$dummy [1450]), .D (nx47270), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47271 (.Y (nx47270), .A0 (ram_107__5), .A1 (nx65650), .S0 (
             nx63740)) ;
    dffr reg_ram_106__5 (.Q (ram_106__5), .QB (\$dummy [1451]), .D (nx47280), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47281 (.Y (nx47280), .A0 (ram_106__5), .A1 (nx65650), .S0 (
             nx63744)) ;
    aoi22 ix60725 (.Y (nx60724), .A0 (ram_108__5), .A1 (nx64970), .B0 (
          ram_109__5), .B1 (nx65008)) ;
    dffr reg_ram_108__5 (.Q (ram_108__5), .QB (\$dummy [1452]), .D (nx47260), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47261 (.Y (nx47260), .A0 (ram_108__5), .A1 (nx65650), .S0 (
             nx63736)) ;
    dffr reg_ram_109__5 (.Q (ram_109__5), .QB (\$dummy [1453]), .D (nx47250), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47251 (.Y (nx47250), .A0 (ram_109__5), .A1 (nx65650), .S0 (
             nx63732)) ;
    aoi22 ix60733 (.Y (nx60732), .A0 (ram_111__5), .A1 (nx65046), .B0 (
          ram_110__5), .B1 (nx65084)) ;
    dffr reg_ram_111__5 (.Q (ram_111__5), .QB (\$dummy [1454]), .D (nx47230), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47231 (.Y (nx47230), .A0 (ram_111__5), .A1 (nx65650), .S0 (
             nx63724)) ;
    dffr reg_ram_110__5 (.Q (ram_110__5), .QB (\$dummy [1455]), .D (nx47240), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47241 (.Y (nx47240), .A0 (ram_110__5), .A1 (nx65652), .S0 (
             nx63728)) ;
    oai21 ix60741 (.Y (nx60740), .A0 (nx16094), .A1 (nx16016), .B0 (nx65210)) ;
    nand04 ix16095 (.Y (nx16094), .A0 (nx60743), .A1 (nx60751), .A2 (nx60759), .A3 (
           nx60767)) ;
    aoi22 ix60744 (.Y (nx60743), .A0 (ram_112__5), .A1 (nx64514), .B0 (
          ram_113__5), .B1 (nx64552)) ;
    dffr reg_ram_112__5 (.Q (ram_112__5), .QB (\$dummy [1456]), .D (nx47220), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47221 (.Y (nx47220), .A0 (ram_112__5), .A1 (nx65652), .S0 (
             nx63714)) ;
    dffr reg_ram_113__5 (.Q (ram_113__5), .QB (\$dummy [1457]), .D (nx47210), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47211 (.Y (nx47210), .A0 (ram_113__5), .A1 (nx65652), .S0 (
             nx63710)) ;
    aoi22 ix60752 (.Y (nx60751), .A0 (ram_115__5), .A1 (nx64590), .B0 (
          ram_114__5), .B1 (nx64628)) ;
    dffr reg_ram_115__5 (.Q (ram_115__5), .QB (\$dummy [1458]), .D (nx47190), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47191 (.Y (nx47190), .A0 (ram_115__5), .A1 (nx65652), .S0 (
             nx63702)) ;
    dffr reg_ram_114__5 (.Q (ram_114__5), .QB (\$dummy [1459]), .D (nx47200), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47201 (.Y (nx47200), .A0 (ram_114__5), .A1 (nx65652), .S0 (
             nx63706)) ;
    aoi22 ix60760 (.Y (nx60759), .A0 (ram_116__5), .A1 (nx64666), .B0 (
          ram_117__5), .B1 (nx64704)) ;
    dffr reg_ram_116__5 (.Q (ram_116__5), .QB (\$dummy [1460]), .D (nx47180), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47181 (.Y (nx47180), .A0 (ram_116__5), .A1 (nx65652), .S0 (
             nx63698)) ;
    dffr reg_ram_117__5 (.Q (ram_117__5), .QB (\$dummy [1461]), .D (nx47170), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47171 (.Y (nx47170), .A0 (ram_117__5), .A1 (nx65652), .S0 (
             nx63694)) ;
    aoi22 ix60768 (.Y (nx60767), .A0 (ram_119__5), .A1 (nx64742), .B0 (
          ram_118__5), .B1 (nx64780)) ;
    dffr reg_ram_119__5 (.Q (ram_119__5), .QB (\$dummy [1462]), .D (nx47150), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47151 (.Y (nx47150), .A0 (ram_119__5), .A1 (nx65654), .S0 (
             nx63686)) ;
    dffr reg_ram_118__5 (.Q (ram_118__5), .QB (\$dummy [1463]), .D (nx47160), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47161 (.Y (nx47160), .A0 (ram_118__5), .A1 (nx65654), .S0 (
             nx63690)) ;
    nand04 ix16017 (.Y (nx16016), .A0 (nx60776), .A1 (nx60784), .A2 (nx60792), .A3 (
           nx60800)) ;
    aoi22 ix60777 (.Y (nx60776), .A0 (ram_120__5), .A1 (nx64818), .B0 (
          ram_121__5), .B1 (nx64856)) ;
    dffr reg_ram_120__5 (.Q (ram_120__5), .QB (\$dummy [1464]), .D (nx47140), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47141 (.Y (nx47140), .A0 (ram_120__5), .A1 (nx65654), .S0 (
             nx63682)) ;
    dffr reg_ram_121__5 (.Q (ram_121__5), .QB (\$dummy [1465]), .D (nx47130), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47131 (.Y (nx47130), .A0 (ram_121__5), .A1 (nx65654), .S0 (
             nx63678)) ;
    aoi22 ix60785 (.Y (nx60784), .A0 (ram_123__5), .A1 (nx64894), .B0 (
          ram_122__5), .B1 (nx64932)) ;
    dffr reg_ram_123__5 (.Q (ram_123__5), .QB (\$dummy [1466]), .D (nx47110), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47111 (.Y (nx47110), .A0 (ram_123__5), .A1 (nx65654), .S0 (
             nx63670)) ;
    dffr reg_ram_122__5 (.Q (ram_122__5), .QB (\$dummy [1467]), .D (nx47120), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47121 (.Y (nx47120), .A0 (ram_122__5), .A1 (nx65654), .S0 (
             nx63674)) ;
    aoi22 ix60793 (.Y (nx60792), .A0 (ram_124__5), .A1 (nx64970), .B0 (
          ram_125__5), .B1 (nx65008)) ;
    dffr reg_ram_124__5 (.Q (ram_124__5), .QB (\$dummy [1468]), .D (nx47100), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47101 (.Y (nx47100), .A0 (ram_124__5), .A1 (nx65654), .S0 (
             nx63666)) ;
    dffr reg_ram_125__5 (.Q (ram_125__5), .QB (\$dummy [1469]), .D (nx47090), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47091 (.Y (nx47090), .A0 (ram_125__5), .A1 (nx65656), .S0 (
             nx63662)) ;
    aoi22 ix60801 (.Y (nx60800), .A0 (ram_127__5), .A1 (nx65046), .B0 (
          ram_126__5), .B1 (nx65084)) ;
    dffr reg_ram_127__5 (.Q (ram_127__5), .QB (\$dummy [1470]), .D (nx47070), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47071 (.Y (nx47070), .A0 (ram_127__5), .A1 (nx65656), .S0 (
             nx63654)) ;
    dffr reg_ram_126__5 (.Q (ram_126__5), .QB (\$dummy [1471]), .D (nx47080), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47081 (.Y (nx47080), .A0 (ram_126__5), .A1 (nx65656), .S0 (
             nx63658)) ;
    nand04 ix15939 (.Y (nx15938), .A0 (nx60809), .A1 (nx60877), .A2 (nx60945), .A3 (
           nx61013)) ;
    oai21 ix60810 (.Y (nx60809), .A0 (nx15928), .A1 (nx15850), .B0 (nx65214)) ;
    nand04 ix15929 (.Y (nx15928), .A0 (nx60812), .A1 (nx60820), .A2 (nx60828), .A3 (
           nx60836)) ;
    aoi22 ix60813 (.Y (nx60812), .A0 (ram_128__5), .A1 (nx64514), .B0 (
          ram_129__5), .B1 (nx64552)) ;
    dffr reg_ram_128__5 (.Q (ram_128__5), .QB (\$dummy [1472]), .D (nx47060), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47061 (.Y (nx47060), .A0 (ram_128__5), .A1 (nx65656), .S0 (
             nx63644)) ;
    dffr reg_ram_129__5 (.Q (ram_129__5), .QB (\$dummy [1473]), .D (nx47050), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47051 (.Y (nx47050), .A0 (ram_129__5), .A1 (nx65656), .S0 (
             nx63640)) ;
    aoi22 ix60821 (.Y (nx60820), .A0 (ram_131__5), .A1 (nx64590), .B0 (
          ram_130__5), .B1 (nx64628)) ;
    dffr reg_ram_131__5 (.Q (ram_131__5), .QB (\$dummy [1474]), .D (nx47030), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47031 (.Y (nx47030), .A0 (ram_131__5), .A1 (nx65656), .S0 (
             nx63632)) ;
    dffr reg_ram_130__5 (.Q (ram_130__5), .QB (\$dummy [1475]), .D (nx47040), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47041 (.Y (nx47040), .A0 (ram_130__5), .A1 (nx65656), .S0 (
             nx63636)) ;
    aoi22 ix60829 (.Y (nx60828), .A0 (ram_132__5), .A1 (nx64666), .B0 (
          ram_133__5), .B1 (nx64704)) ;
    dffr reg_ram_132__5 (.Q (ram_132__5), .QB (\$dummy [1476]), .D (nx47020), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47021 (.Y (nx47020), .A0 (ram_132__5), .A1 (nx65658), .S0 (
             nx63628)) ;
    dffr reg_ram_133__5 (.Q (ram_133__5), .QB (\$dummy [1477]), .D (nx47010), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47011 (.Y (nx47010), .A0 (ram_133__5), .A1 (nx65658), .S0 (
             nx63624)) ;
    aoi22 ix60837 (.Y (nx60836), .A0 (ram_135__5), .A1 (nx64742), .B0 (
          ram_134__5), .B1 (nx64780)) ;
    dffr reg_ram_135__5 (.Q (ram_135__5), .QB (\$dummy [1478]), .D (nx46990), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46991 (.Y (nx46990), .A0 (ram_135__5), .A1 (nx65658), .S0 (
             nx63616)) ;
    dffr reg_ram_134__5 (.Q (ram_134__5), .QB (\$dummy [1479]), .D (nx47000), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix47001 (.Y (nx47000), .A0 (ram_134__5), .A1 (nx65658), .S0 (
             nx63620)) ;
    nand04 ix15851 (.Y (nx15850), .A0 (nx60845), .A1 (nx60853), .A2 (nx60861), .A3 (
           nx60869)) ;
    aoi22 ix60846 (.Y (nx60845), .A0 (ram_136__5), .A1 (nx64818), .B0 (
          ram_137__5), .B1 (nx64856)) ;
    dffr reg_ram_136__5 (.Q (ram_136__5), .QB (\$dummy [1480]), .D (nx46980), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46981 (.Y (nx46980), .A0 (ram_136__5), .A1 (nx65658), .S0 (
             nx63612)) ;
    dffr reg_ram_137__5 (.Q (ram_137__5), .QB (\$dummy [1481]), .D (nx46970), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46971 (.Y (nx46970), .A0 (ram_137__5), .A1 (nx65658), .S0 (
             nx63608)) ;
    aoi22 ix60854 (.Y (nx60853), .A0 (ram_139__5), .A1 (nx64894), .B0 (
          ram_138__5), .B1 (nx64932)) ;
    dffr reg_ram_139__5 (.Q (ram_139__5), .QB (\$dummy [1482]), .D (nx46950), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46951 (.Y (nx46950), .A0 (ram_139__5), .A1 (nx65658), .S0 (
             nx63600)) ;
    dffr reg_ram_138__5 (.Q (ram_138__5), .QB (\$dummy [1483]), .D (nx46960), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46961 (.Y (nx46960), .A0 (ram_138__5), .A1 (nx65660), .S0 (
             nx63604)) ;
    aoi22 ix60862 (.Y (nx60861), .A0 (ram_140__5), .A1 (nx64970), .B0 (
          ram_141__5), .B1 (nx65008)) ;
    dffr reg_ram_140__5 (.Q (ram_140__5), .QB (\$dummy [1484]), .D (nx46940), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46941 (.Y (nx46940), .A0 (ram_140__5), .A1 (nx65660), .S0 (
             nx63596)) ;
    dffr reg_ram_141__5 (.Q (ram_141__5), .QB (\$dummy [1485]), .D (nx46930), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46931 (.Y (nx46930), .A0 (ram_141__5), .A1 (nx65660), .S0 (
             nx63592)) ;
    aoi22 ix60870 (.Y (nx60869), .A0 (ram_143__5), .A1 (nx65046), .B0 (
          ram_142__5), .B1 (nx65084)) ;
    dffr reg_ram_143__5 (.Q (ram_143__5), .QB (\$dummy [1486]), .D (nx46910), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46911 (.Y (nx46910), .A0 (ram_143__5), .A1 (nx65660), .S0 (
             nx63584)) ;
    dffr reg_ram_142__5 (.Q (ram_142__5), .QB (\$dummy [1487]), .D (nx46920), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46921 (.Y (nx46920), .A0 (ram_142__5), .A1 (nx65660), .S0 (
             nx63588)) ;
    oai21 ix60878 (.Y (nx60877), .A0 (nx15766), .A1 (nx15688), .B0 (nx65218)) ;
    nand04 ix15767 (.Y (nx15766), .A0 (nx60880), .A1 (nx60888), .A2 (nx60896), .A3 (
           nx60904)) ;
    aoi22 ix60881 (.Y (nx60880), .A0 (ram_144__5), .A1 (nx64514), .B0 (
          ram_145__5), .B1 (nx64552)) ;
    dffr reg_ram_144__5 (.Q (ram_144__5), .QB (\$dummy [1488]), .D (nx46900), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46901 (.Y (nx46900), .A0 (ram_144__5), .A1 (nx65660), .S0 (
             nx63574)) ;
    dffr reg_ram_145__5 (.Q (ram_145__5), .QB (\$dummy [1489]), .D (nx46890), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46891 (.Y (nx46890), .A0 (ram_145__5), .A1 (nx65660), .S0 (
             nx63570)) ;
    aoi22 ix60889 (.Y (nx60888), .A0 (ram_147__5), .A1 (nx64590), .B0 (
          ram_146__5), .B1 (nx64628)) ;
    dffr reg_ram_147__5 (.Q (ram_147__5), .QB (\$dummy [1490]), .D (nx46870), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46871 (.Y (nx46870), .A0 (ram_147__5), .A1 (nx65662), .S0 (
             nx63562)) ;
    dffr reg_ram_146__5 (.Q (ram_146__5), .QB (\$dummy [1491]), .D (nx46880), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46881 (.Y (nx46880), .A0 (ram_146__5), .A1 (nx65662), .S0 (
             nx63566)) ;
    aoi22 ix60897 (.Y (nx60896), .A0 (ram_148__5), .A1 (nx64666), .B0 (
          ram_149__5), .B1 (nx64704)) ;
    dffr reg_ram_148__5 (.Q (ram_148__5), .QB (\$dummy [1492]), .D (nx46860), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46861 (.Y (nx46860), .A0 (ram_148__5), .A1 (nx65662), .S0 (
             nx63558)) ;
    dffr reg_ram_149__5 (.Q (ram_149__5), .QB (\$dummy [1493]), .D (nx46850), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46851 (.Y (nx46850), .A0 (ram_149__5), .A1 (nx65662), .S0 (
             nx63554)) ;
    aoi22 ix60905 (.Y (nx60904), .A0 (ram_151__5), .A1 (nx64742), .B0 (
          ram_150__5), .B1 (nx64780)) ;
    dffr reg_ram_151__5 (.Q (ram_151__5), .QB (\$dummy [1494]), .D (nx46830), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46831 (.Y (nx46830), .A0 (ram_151__5), .A1 (nx65662), .S0 (
             nx63546)) ;
    dffr reg_ram_150__5 (.Q (ram_150__5), .QB (\$dummy [1495]), .D (nx46840), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46841 (.Y (nx46840), .A0 (ram_150__5), .A1 (nx65662), .S0 (
             nx63550)) ;
    nand04 ix15689 (.Y (nx15688), .A0 (nx60913), .A1 (nx60921), .A2 (nx60929), .A3 (
           nx60937)) ;
    aoi22 ix60914 (.Y (nx60913), .A0 (ram_152__5), .A1 (nx64818), .B0 (
          ram_153__5), .B1 (nx64856)) ;
    dffr reg_ram_152__5 (.Q (ram_152__5), .QB (\$dummy [1496]), .D (nx46820), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46821 (.Y (nx46820), .A0 (ram_152__5), .A1 (nx65662), .S0 (
             nx63542)) ;
    dffr reg_ram_153__5 (.Q (ram_153__5), .QB (\$dummy [1497]), .D (nx46810), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46811 (.Y (nx46810), .A0 (ram_153__5), .A1 (nx65664), .S0 (
             nx63538)) ;
    aoi22 ix60922 (.Y (nx60921), .A0 (ram_155__5), .A1 (nx64894), .B0 (
          ram_154__5), .B1 (nx64932)) ;
    dffr reg_ram_155__5 (.Q (ram_155__5), .QB (\$dummy [1498]), .D (nx46790), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46791 (.Y (nx46790), .A0 (ram_155__5), .A1 (nx65664), .S0 (
             nx63530)) ;
    dffr reg_ram_154__5 (.Q (ram_154__5), .QB (\$dummy [1499]), .D (nx46800), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46801 (.Y (nx46800), .A0 (ram_154__5), .A1 (nx65664), .S0 (
             nx63534)) ;
    aoi22 ix60930 (.Y (nx60929), .A0 (ram_156__5), .A1 (nx64970), .B0 (
          ram_157__5), .B1 (nx65008)) ;
    dffr reg_ram_156__5 (.Q (ram_156__5), .QB (\$dummy [1500]), .D (nx46780), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46781 (.Y (nx46780), .A0 (ram_156__5), .A1 (nx65664), .S0 (
             nx63526)) ;
    dffr reg_ram_157__5 (.Q (ram_157__5), .QB (\$dummy [1501]), .D (nx46770), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46771 (.Y (nx46770), .A0 (ram_157__5), .A1 (nx65664), .S0 (
             nx63522)) ;
    aoi22 ix60938 (.Y (nx60937), .A0 (ram_159__5), .A1 (nx65046), .B0 (
          ram_158__5), .B1 (nx65084)) ;
    dffr reg_ram_159__5 (.Q (ram_159__5), .QB (\$dummy [1502]), .D (nx46750), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46751 (.Y (nx46750), .A0 (ram_159__5), .A1 (nx65664), .S0 (
             nx63514)) ;
    dffr reg_ram_158__5 (.Q (ram_158__5), .QB (\$dummy [1503]), .D (nx46760), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46761 (.Y (nx46760), .A0 (ram_158__5), .A1 (nx65664), .S0 (
             nx63518)) ;
    oai21 ix60946 (.Y (nx60945), .A0 (nx15602), .A1 (nx15524), .B0 (nx65222)) ;
    nand04 ix15603 (.Y (nx15602), .A0 (nx60948), .A1 (nx60956), .A2 (nx60964), .A3 (
           nx60972)) ;
    aoi22 ix60949 (.Y (nx60948), .A0 (ram_160__5), .A1 (nx64514), .B0 (
          ram_161__5), .B1 (nx64552)) ;
    dffr reg_ram_160__5 (.Q (ram_160__5), .QB (\$dummy [1504]), .D (nx46740), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46741 (.Y (nx46740), .A0 (ram_160__5), .A1 (nx65666), .S0 (
             nx63504)) ;
    dffr reg_ram_161__5 (.Q (ram_161__5), .QB (\$dummy [1505]), .D (nx46730), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46731 (.Y (nx46730), .A0 (ram_161__5), .A1 (nx65666), .S0 (
             nx63500)) ;
    aoi22 ix60957 (.Y (nx60956), .A0 (ram_163__5), .A1 (nx64590), .B0 (
          ram_162__5), .B1 (nx64628)) ;
    dffr reg_ram_163__5 (.Q (ram_163__5), .QB (\$dummy [1506]), .D (nx46710), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46711 (.Y (nx46710), .A0 (ram_163__5), .A1 (nx65666), .S0 (
             nx63492)) ;
    dffr reg_ram_162__5 (.Q (ram_162__5), .QB (\$dummy [1507]), .D (nx46720), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46721 (.Y (nx46720), .A0 (ram_162__5), .A1 (nx65666), .S0 (
             nx63496)) ;
    aoi22 ix60965 (.Y (nx60964), .A0 (ram_164__5), .A1 (nx64666), .B0 (
          ram_165__5), .B1 (nx64704)) ;
    dffr reg_ram_164__5 (.Q (ram_164__5), .QB (\$dummy [1508]), .D (nx46700), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46701 (.Y (nx46700), .A0 (ram_164__5), .A1 (nx65666), .S0 (
             nx63488)) ;
    dffr reg_ram_165__5 (.Q (ram_165__5), .QB (\$dummy [1509]), .D (nx46690), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46691 (.Y (nx46690), .A0 (ram_165__5), .A1 (nx65666), .S0 (
             nx63484)) ;
    aoi22 ix60973 (.Y (nx60972), .A0 (ram_167__5), .A1 (nx64742), .B0 (
          ram_166__5), .B1 (nx64780)) ;
    dffr reg_ram_167__5 (.Q (ram_167__5), .QB (\$dummy [1510]), .D (nx46670), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46671 (.Y (nx46670), .A0 (ram_167__5), .A1 (nx65666), .S0 (
             nx63476)) ;
    dffr reg_ram_166__5 (.Q (ram_166__5), .QB (\$dummy [1511]), .D (nx46680), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46681 (.Y (nx46680), .A0 (ram_166__5), .A1 (nx65668), .S0 (
             nx63480)) ;
    nand04 ix15525 (.Y (nx15524), .A0 (nx60981), .A1 (nx60989), .A2 (nx60997), .A3 (
           nx61005)) ;
    aoi22 ix60982 (.Y (nx60981), .A0 (ram_168__5), .A1 (nx64818), .B0 (
          ram_169__5), .B1 (nx64856)) ;
    dffr reg_ram_168__5 (.Q (ram_168__5), .QB (\$dummy [1512]), .D (nx46660), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46661 (.Y (nx46660), .A0 (ram_168__5), .A1 (nx65668), .S0 (
             nx63472)) ;
    dffr reg_ram_169__5 (.Q (ram_169__5), .QB (\$dummy [1513]), .D (nx46650), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46651 (.Y (nx46650), .A0 (ram_169__5), .A1 (nx65668), .S0 (
             nx63468)) ;
    aoi22 ix60990 (.Y (nx60989), .A0 (ram_171__5), .A1 (nx64894), .B0 (
          ram_170__5), .B1 (nx64932)) ;
    dffr reg_ram_171__5 (.Q (ram_171__5), .QB (\$dummy [1514]), .D (nx46630), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46631 (.Y (nx46630), .A0 (ram_171__5), .A1 (nx65668), .S0 (
             nx63460)) ;
    dffr reg_ram_170__5 (.Q (ram_170__5), .QB (\$dummy [1515]), .D (nx46640), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46641 (.Y (nx46640), .A0 (ram_170__5), .A1 (nx65668), .S0 (
             nx63464)) ;
    aoi22 ix60998 (.Y (nx60997), .A0 (ram_172__5), .A1 (nx64970), .B0 (
          ram_173__5), .B1 (nx65008)) ;
    dffr reg_ram_172__5 (.Q (ram_172__5), .QB (\$dummy [1516]), .D (nx46620), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46621 (.Y (nx46620), .A0 (ram_172__5), .A1 (nx65668), .S0 (
             nx63456)) ;
    dffr reg_ram_173__5 (.Q (ram_173__5), .QB (\$dummy [1517]), .D (nx46610), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46611 (.Y (nx46610), .A0 (ram_173__5), .A1 (nx65668), .S0 (
             nx63452)) ;
    aoi22 ix61006 (.Y (nx61005), .A0 (ram_175__5), .A1 (nx65046), .B0 (
          ram_174__5), .B1 (nx65084)) ;
    dffr reg_ram_175__5 (.Q (ram_175__5), .QB (\$dummy [1518]), .D (nx46590), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46591 (.Y (nx46590), .A0 (ram_175__5), .A1 (nx65670), .S0 (
             nx63444)) ;
    dffr reg_ram_174__5 (.Q (ram_174__5), .QB (\$dummy [1519]), .D (nx46600), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46601 (.Y (nx46600), .A0 (ram_174__5), .A1 (nx65670), .S0 (
             nx63448)) ;
    oai21 ix61014 (.Y (nx61013), .A0 (nx15440), .A1 (nx15362), .B0 (nx65226)) ;
    nand04 ix15441 (.Y (nx15440), .A0 (nx61016), .A1 (nx61024), .A2 (nx61032), .A3 (
           nx61040)) ;
    aoi22 ix61017 (.Y (nx61016), .A0 (ram_176__5), .A1 (nx64514), .B0 (
          ram_177__5), .B1 (nx64552)) ;
    dffr reg_ram_176__5 (.Q (ram_176__5), .QB (\$dummy [1520]), .D (nx46580), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46581 (.Y (nx46580), .A0 (ram_176__5), .A1 (nx65670), .S0 (
             nx63434)) ;
    dffr reg_ram_177__5 (.Q (ram_177__5), .QB (\$dummy [1521]), .D (nx46570), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46571 (.Y (nx46570), .A0 (ram_177__5), .A1 (nx65670), .S0 (
             nx63424)) ;
    aoi22 ix61025 (.Y (nx61024), .A0 (ram_179__5), .A1 (nx64590), .B0 (
          ram_178__5), .B1 (nx64628)) ;
    dffr reg_ram_179__5 (.Q (ram_179__5), .QB (\$dummy [1522]), .D (nx46550), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46551 (.Y (nx46550), .A0 (ram_179__5), .A1 (nx65670), .S0 (
             nx63404)) ;
    dffr reg_ram_178__5 (.Q (ram_178__5), .QB (\$dummy [1523]), .D (nx46560), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46561 (.Y (nx46560), .A0 (ram_178__5), .A1 (nx65670), .S0 (
             nx63414)) ;
    aoi22 ix61033 (.Y (nx61032), .A0 (ram_180__5), .A1 (nx64666), .B0 (
          ram_181__5), .B1 (nx64704)) ;
    dffr reg_ram_180__5 (.Q (ram_180__5), .QB (\$dummy [1524]), .D (nx46540), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46541 (.Y (nx46540), .A0 (ram_180__5), .A1 (nx65670), .S0 (
             nx63394)) ;
    dffr reg_ram_181__5 (.Q (ram_181__5), .QB (\$dummy [1525]), .D (nx46530), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46531 (.Y (nx46530), .A0 (ram_181__5), .A1 (nx65672), .S0 (
             nx63384)) ;
    aoi22 ix61041 (.Y (nx61040), .A0 (ram_183__5), .A1 (nx64742), .B0 (
          ram_182__5), .B1 (nx64780)) ;
    dffr reg_ram_183__5 (.Q (ram_183__5), .QB (\$dummy [1526]), .D (nx46510), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46511 (.Y (nx46510), .A0 (ram_183__5), .A1 (nx65672), .S0 (
             nx63364)) ;
    dffr reg_ram_182__5 (.Q (ram_182__5), .QB (\$dummy [1527]), .D (nx46520), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46521 (.Y (nx46520), .A0 (ram_182__5), .A1 (nx65672), .S0 (
             nx63374)) ;
    nand04 ix15363 (.Y (nx15362), .A0 (nx61049), .A1 (nx61057), .A2 (nx61065), .A3 (
           nx61073)) ;
    aoi22 ix61050 (.Y (nx61049), .A0 (ram_184__5), .A1 (nx64818), .B0 (
          ram_185__5), .B1 (nx64856)) ;
    dffr reg_ram_184__5 (.Q (ram_184__5), .QB (\$dummy [1528]), .D (nx46500), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46501 (.Y (nx46500), .A0 (ram_184__5), .A1 (nx65672), .S0 (
             nx63354)) ;
    dffr reg_ram_185__5 (.Q (ram_185__5), .QB (\$dummy [1529]), .D (nx46490), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46491 (.Y (nx46490), .A0 (ram_185__5), .A1 (nx65672), .S0 (
             nx63344)) ;
    aoi22 ix61058 (.Y (nx61057), .A0 (ram_187__5), .A1 (nx64894), .B0 (
          ram_186__5), .B1 (nx64932)) ;
    dffr reg_ram_187__5 (.Q (ram_187__5), .QB (\$dummy [1530]), .D (nx46470), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46471 (.Y (nx46470), .A0 (ram_187__5), .A1 (nx65672), .S0 (
             nx63324)) ;
    dffr reg_ram_186__5 (.Q (ram_186__5), .QB (\$dummy [1531]), .D (nx46480), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46481 (.Y (nx46480), .A0 (ram_186__5), .A1 (nx65672), .S0 (
             nx63334)) ;
    aoi22 ix61066 (.Y (nx61065), .A0 (ram_188__5), .A1 (nx64970), .B0 (
          ram_189__5), .B1 (nx65008)) ;
    dffr reg_ram_188__5 (.Q (ram_188__5), .QB (\$dummy [1532]), .D (nx46460), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46461 (.Y (nx46460), .A0 (ram_188__5), .A1 (nx65674), .S0 (
             nx63314)) ;
    dffr reg_ram_189__5 (.Q (ram_189__5), .QB (\$dummy [1533]), .D (nx46450), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46451 (.Y (nx46450), .A0 (ram_189__5), .A1 (nx65674), .S0 (
             nx63304)) ;
    aoi22 ix61074 (.Y (nx61073), .A0 (ram_191__5), .A1 (nx65046), .B0 (
          ram_190__5), .B1 (nx65084)) ;
    dffr reg_ram_191__5 (.Q (ram_191__5), .QB (\$dummy [1534]), .D (nx46430), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46431 (.Y (nx46430), .A0 (ram_191__5), .A1 (nx65674), .S0 (
             nx63284)) ;
    dffr reg_ram_190__5 (.Q (ram_190__5), .QB (\$dummy [1535]), .D (nx46440), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix46441 (.Y (nx46440), .A0 (ram_190__5), .A1 (nx65674), .S0 (
             nx63294)) ;
    or04 ix20529 (.Y (dataout[6]), .A0 (nx20524), .A1 (nx19870), .A2 (nx19214), 
         .A3 (nx18560)) ;
    nand04 ix20525 (.Y (nx20524), .A0 (nx61083), .A1 (nx61151), .A2 (nx61219), .A3 (
           nx61287)) ;
    oai21 ix61084 (.Y (nx61083), .A0 (nx20514), .A1 (nx20436), .B0 (nx65096)) ;
    nand04 ix20515 (.Y (nx20514), .A0 (nx61086), .A1 (nx61094), .A2 (nx61102), .A3 (
           nx61110)) ;
    aoi22 ix61087 (.Y (nx61086), .A0 (ram_240__6), .A1 (nx64514), .B0 (
          ram_241__6), .B1 (nx64552)) ;
    dffr reg_ram_240__6 (.Q (ram_240__6), .QB (\$dummy [1536]), .D (nx51540), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51541 (.Y (nx51540), .A0 (ram_240__6), .A1 (nx65526), .S0 (
             nx64414)) ;
    dffr reg_ram_241__6 (.Q (ram_241__6), .QB (\$dummy [1537]), .D (nx51530), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51531 (.Y (nx51530), .A0 (ram_241__6), .A1 (nx65526), .S0 (
             nx64410)) ;
    aoi22 ix61095 (.Y (nx61094), .A0 (ram_243__6), .A1 (nx64590), .B0 (
          ram_242__6), .B1 (nx64628)) ;
    dffr reg_ram_243__6 (.Q (ram_243__6), .QB (\$dummy [1538]), .D (nx51510), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51511 (.Y (nx51510), .A0 (ram_243__6), .A1 (nx65526), .S0 (
             nx64402)) ;
    dffr reg_ram_242__6 (.Q (ram_242__6), .QB (\$dummy [1539]), .D (nx51520), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51521 (.Y (nx51520), .A0 (ram_242__6), .A1 (nx65526), .S0 (
             nx64406)) ;
    aoi22 ix61103 (.Y (nx61102), .A0 (ram_244__6), .A1 (nx64666), .B0 (
          ram_245__6), .B1 (nx64704)) ;
    dffr reg_ram_244__6 (.Q (ram_244__6), .QB (\$dummy [1540]), .D (nx51500), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51501 (.Y (nx51500), .A0 (ram_244__6), .A1 (nx65526), .S0 (
             nx64398)) ;
    dffr reg_ram_245__6 (.Q (ram_245__6), .QB (\$dummy [1541]), .D (nx51490), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51491 (.Y (nx51490), .A0 (ram_245__6), .A1 (nx65526), .S0 (
             nx64394)) ;
    aoi22 ix61111 (.Y (nx61110), .A0 (ram_247__6), .A1 (nx64742), .B0 (
          ram_246__6), .B1 (nx64780)) ;
    dffr reg_ram_247__6 (.Q (ram_247__6), .QB (\$dummy [1542]), .D (nx51470), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51471 (.Y (nx51470), .A0 (ram_247__6), .A1 (nx65526), .S0 (
             nx64386)) ;
    dffr reg_ram_246__6 (.Q (ram_246__6), .QB (\$dummy [1543]), .D (nx51480), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51481 (.Y (nx51480), .A0 (ram_246__6), .A1 (nx65528), .S0 (
             nx64390)) ;
    nand04 ix20437 (.Y (nx20436), .A0 (nx61119), .A1 (nx61127), .A2 (nx61135), .A3 (
           nx61143)) ;
    aoi22 ix61120 (.Y (nx61119), .A0 (ram_248__6), .A1 (nx64818), .B0 (
          ram_249__6), .B1 (nx64856)) ;
    dffr reg_ram_248__6 (.Q (ram_248__6), .QB (\$dummy [1544]), .D (nx51460), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51461 (.Y (nx51460), .A0 (ram_248__6), .A1 (nx65528), .S0 (
             nx64382)) ;
    dffr reg_ram_249__6 (.Q (ram_249__6), .QB (\$dummy [1545]), .D (nx51450), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51451 (.Y (nx51450), .A0 (ram_249__6), .A1 (nx65528), .S0 (
             nx64378)) ;
    aoi22 ix61128 (.Y (nx61127), .A0 (ram_251__6), .A1 (nx64894), .B0 (
          ram_250__6), .B1 (nx64932)) ;
    dffr reg_ram_251__6 (.Q (ram_251__6), .QB (\$dummy [1546]), .D (nx51430), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51431 (.Y (nx51430), .A0 (ram_251__6), .A1 (nx65528), .S0 (
             nx64370)) ;
    dffr reg_ram_250__6 (.Q (ram_250__6), .QB (\$dummy [1547]), .D (nx51440), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51441 (.Y (nx51440), .A0 (ram_250__6), .A1 (nx65528), .S0 (
             nx64374)) ;
    aoi22 ix61136 (.Y (nx61135), .A0 (ram_252__6), .A1 (nx64970), .B0 (
          ram_253__6), .B1 (nx65008)) ;
    dffr reg_ram_252__6 (.Q (ram_252__6), .QB (\$dummy [1548]), .D (nx51420), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51421 (.Y (nx51420), .A0 (ram_252__6), .A1 (nx65528), .S0 (
             nx64366)) ;
    dffr reg_ram_253__6 (.Q (ram_253__6), .QB (\$dummy [1549]), .D (nx51410), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51411 (.Y (nx51410), .A0 (ram_253__6), .A1 (nx65528), .S0 (
             nx64362)) ;
    aoi22 ix61144 (.Y (nx61143), .A0 (ram_255__6), .A1 (nx65046), .B0 (
          ram_254__6), .B1 (nx65084)) ;
    dffr reg_ram_255__6 (.Q (ram_255__6), .QB (\$dummy [1550]), .D (nx51390), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51391 (.Y (nx51390), .A0 (ram_255__6), .A1 (nx65530), .S0 (
             nx64354)) ;
    dffr reg_ram_254__6 (.Q (ram_254__6), .QB (\$dummy [1551]), .D (nx51400), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51401 (.Y (nx51400), .A0 (ram_254__6), .A1 (nx65530), .S0 (
             nx64358)) ;
    oai21 ix61152 (.Y (nx61151), .A0 (nx20352), .A1 (nx20274), .B0 (nx65100)) ;
    nand04 ix20353 (.Y (nx20352), .A0 (nx61154), .A1 (nx61162), .A2 (nx61170), .A3 (
           nx61178)) ;
    aoi22 ix61155 (.Y (nx61154), .A0 (ram_224__6), .A1 (nx64516), .B0 (
          ram_225__6), .B1 (nx64554)) ;
    dffr reg_ram_224__6 (.Q (ram_224__6), .QB (\$dummy [1552]), .D (nx51380), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51381 (.Y (nx51380), .A0 (ram_224__6), .A1 (nx65530), .S0 (
             nx64344)) ;
    dffr reg_ram_225__6 (.Q (ram_225__6), .QB (\$dummy [1553]), .D (nx51370), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51371 (.Y (nx51370), .A0 (ram_225__6), .A1 (nx65530), .S0 (
             nx64340)) ;
    aoi22 ix61163 (.Y (nx61162), .A0 (ram_227__6), .A1 (nx64592), .B0 (
          ram_226__6), .B1 (nx64630)) ;
    dffr reg_ram_227__6 (.Q (ram_227__6), .QB (\$dummy [1554]), .D (nx51350), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51351 (.Y (nx51350), .A0 (ram_227__6), .A1 (nx65530), .S0 (
             nx64332)) ;
    dffr reg_ram_226__6 (.Q (ram_226__6), .QB (\$dummy [1555]), .D (nx51360), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51361 (.Y (nx51360), .A0 (ram_226__6), .A1 (nx65530), .S0 (
             nx64336)) ;
    aoi22 ix61171 (.Y (nx61170), .A0 (ram_228__6), .A1 (nx64668), .B0 (
          ram_229__6), .B1 (nx64706)) ;
    dffr reg_ram_228__6 (.Q (ram_228__6), .QB (\$dummy [1556]), .D (nx51340), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51341 (.Y (nx51340), .A0 (ram_228__6), .A1 (nx65530), .S0 (
             nx64328)) ;
    dffr reg_ram_229__6 (.Q (ram_229__6), .QB (\$dummy [1557]), .D (nx51330), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51331 (.Y (nx51330), .A0 (ram_229__6), .A1 (nx65532), .S0 (
             nx64324)) ;
    aoi22 ix61179 (.Y (nx61178), .A0 (ram_231__6), .A1 (nx64744), .B0 (
          ram_230__6), .B1 (nx64782)) ;
    dffr reg_ram_231__6 (.Q (ram_231__6), .QB (\$dummy [1558]), .D (nx51310), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51311 (.Y (nx51310), .A0 (ram_231__6), .A1 (nx65532), .S0 (
             nx64316)) ;
    dffr reg_ram_230__6 (.Q (ram_230__6), .QB (\$dummy [1559]), .D (nx51320), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51321 (.Y (nx51320), .A0 (ram_230__6), .A1 (nx65532), .S0 (
             nx64320)) ;
    nand04 ix20275 (.Y (nx20274), .A0 (nx61187), .A1 (nx61195), .A2 (nx61203), .A3 (
           nx61211)) ;
    aoi22 ix61188 (.Y (nx61187), .A0 (ram_232__6), .A1 (nx64820), .B0 (
          ram_233__6), .B1 (nx64858)) ;
    dffr reg_ram_232__6 (.Q (ram_232__6), .QB (\$dummy [1560]), .D (nx51300), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51301 (.Y (nx51300), .A0 (ram_232__6), .A1 (nx65532), .S0 (
             nx64312)) ;
    dffr reg_ram_233__6 (.Q (ram_233__6), .QB (\$dummy [1561]), .D (nx51290), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51291 (.Y (nx51290), .A0 (ram_233__6), .A1 (nx65532), .S0 (
             nx64308)) ;
    aoi22 ix61196 (.Y (nx61195), .A0 (ram_235__6), .A1 (nx64896), .B0 (
          ram_234__6), .B1 (nx64934)) ;
    dffr reg_ram_235__6 (.Q (ram_235__6), .QB (\$dummy [1562]), .D (nx51270), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51271 (.Y (nx51270), .A0 (ram_235__6), .A1 (nx65532), .S0 (
             nx64300)) ;
    dffr reg_ram_234__6 (.Q (ram_234__6), .QB (\$dummy [1563]), .D (nx51280), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51281 (.Y (nx51280), .A0 (ram_234__6), .A1 (nx65532), .S0 (
             nx64304)) ;
    aoi22 ix61204 (.Y (nx61203), .A0 (ram_236__6), .A1 (nx64972), .B0 (
          ram_237__6), .B1 (nx65010)) ;
    dffr reg_ram_236__6 (.Q (ram_236__6), .QB (\$dummy [1564]), .D (nx51260), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51261 (.Y (nx51260), .A0 (ram_236__6), .A1 (nx65534), .S0 (
             nx64296)) ;
    dffr reg_ram_237__6 (.Q (ram_237__6), .QB (\$dummy [1565]), .D (nx51250), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51251 (.Y (nx51250), .A0 (ram_237__6), .A1 (nx65534), .S0 (
             nx64292)) ;
    aoi22 ix61212 (.Y (nx61211), .A0 (ram_239__6), .A1 (nx65048), .B0 (
          ram_238__6), .B1 (nx65086)) ;
    dffr reg_ram_239__6 (.Q (ram_239__6), .QB (\$dummy [1566]), .D (nx51230), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51231 (.Y (nx51230), .A0 (ram_239__6), .A1 (nx65534), .S0 (
             nx64284)) ;
    dffr reg_ram_238__6 (.Q (ram_238__6), .QB (\$dummy [1567]), .D (nx51240), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51241 (.Y (nx51240), .A0 (ram_238__6), .A1 (nx65534), .S0 (
             nx64288)) ;
    oai21 ix61220 (.Y (nx61219), .A0 (nx20188), .A1 (nx20110), .B0 (nx65104)) ;
    nand04 ix20189 (.Y (nx20188), .A0 (nx61222), .A1 (nx61230), .A2 (nx61238), .A3 (
           nx61246)) ;
    aoi22 ix61223 (.Y (nx61222), .A0 (ram_208__6), .A1 (nx64516), .B0 (
          ram_209__6), .B1 (nx64554)) ;
    dffr reg_ram_208__6 (.Q (ram_208__6), .QB (\$dummy [1568]), .D (nx51220), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51221 (.Y (nx51220), .A0 (ram_208__6), .A1 (nx65534), .S0 (
             nx64274)) ;
    dffr reg_ram_209__6 (.Q (ram_209__6), .QB (\$dummy [1569]), .D (nx51210), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51211 (.Y (nx51210), .A0 (ram_209__6), .A1 (nx65534), .S0 (
             nx64270)) ;
    aoi22 ix61231 (.Y (nx61230), .A0 (ram_211__6), .A1 (nx64592), .B0 (
          ram_210__6), .B1 (nx64630)) ;
    dffr reg_ram_211__6 (.Q (ram_211__6), .QB (\$dummy [1570]), .D (nx51190), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51191 (.Y (nx51190), .A0 (ram_211__6), .A1 (nx65534), .S0 (
             nx64262)) ;
    dffr reg_ram_210__6 (.Q (ram_210__6), .QB (\$dummy [1571]), .D (nx51200), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51201 (.Y (nx51200), .A0 (ram_210__6), .A1 (nx65536), .S0 (
             nx64266)) ;
    aoi22 ix61239 (.Y (nx61238), .A0 (ram_212__6), .A1 (nx64668), .B0 (
          ram_213__6), .B1 (nx64706)) ;
    dffr reg_ram_212__6 (.Q (ram_212__6), .QB (\$dummy [1572]), .D (nx51180), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51181 (.Y (nx51180), .A0 (ram_212__6), .A1 (nx65536), .S0 (
             nx64258)) ;
    dffr reg_ram_213__6 (.Q (ram_213__6), .QB (\$dummy [1573]), .D (nx51170), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51171 (.Y (nx51170), .A0 (ram_213__6), .A1 (nx65536), .S0 (
             nx64254)) ;
    aoi22 ix61247 (.Y (nx61246), .A0 (ram_215__6), .A1 (nx64744), .B0 (
          ram_214__6), .B1 (nx64782)) ;
    dffr reg_ram_215__6 (.Q (ram_215__6), .QB (\$dummy [1574]), .D (nx51150), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51151 (.Y (nx51150), .A0 (ram_215__6), .A1 (nx65536), .S0 (
             nx64246)) ;
    dffr reg_ram_214__6 (.Q (ram_214__6), .QB (\$dummy [1575]), .D (nx51160), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51161 (.Y (nx51160), .A0 (ram_214__6), .A1 (nx65536), .S0 (
             nx64250)) ;
    nand04 ix20111 (.Y (nx20110), .A0 (nx61255), .A1 (nx61263), .A2 (nx61271), .A3 (
           nx61279)) ;
    aoi22 ix61256 (.Y (nx61255), .A0 (ram_216__6), .A1 (nx64820), .B0 (
          ram_217__6), .B1 (nx64858)) ;
    dffr reg_ram_216__6 (.Q (ram_216__6), .QB (\$dummy [1576]), .D (nx51140), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51141 (.Y (nx51140), .A0 (ram_216__6), .A1 (nx65536), .S0 (
             nx64242)) ;
    dffr reg_ram_217__6 (.Q (ram_217__6), .QB (\$dummy [1577]), .D (nx51130), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51131 (.Y (nx51130), .A0 (ram_217__6), .A1 (nx65536), .S0 (
             nx64238)) ;
    aoi22 ix61264 (.Y (nx61263), .A0 (ram_219__6), .A1 (nx64896), .B0 (
          ram_218__6), .B1 (nx64934)) ;
    dffr reg_ram_219__6 (.Q (ram_219__6), .QB (\$dummy [1578]), .D (nx51110), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51111 (.Y (nx51110), .A0 (ram_219__6), .A1 (nx65538), .S0 (
             nx64230)) ;
    dffr reg_ram_218__6 (.Q (ram_218__6), .QB (\$dummy [1579]), .D (nx51120), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51121 (.Y (nx51120), .A0 (ram_218__6), .A1 (nx65538), .S0 (
             nx64234)) ;
    aoi22 ix61272 (.Y (nx61271), .A0 (ram_220__6), .A1 (nx64972), .B0 (
          ram_221__6), .B1 (nx65010)) ;
    dffr reg_ram_220__6 (.Q (ram_220__6), .QB (\$dummy [1580]), .D (nx51100), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51101 (.Y (nx51100), .A0 (ram_220__6), .A1 (nx65538), .S0 (
             nx64226)) ;
    dffr reg_ram_221__6 (.Q (ram_221__6), .QB (\$dummy [1581]), .D (nx51090), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51091 (.Y (nx51090), .A0 (ram_221__6), .A1 (nx65538), .S0 (
             nx64222)) ;
    aoi22 ix61280 (.Y (nx61279), .A0 (ram_223__6), .A1 (nx65048), .B0 (
          ram_222__6), .B1 (nx65086)) ;
    dffr reg_ram_223__6 (.Q (ram_223__6), .QB (\$dummy [1582]), .D (nx51070), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51071 (.Y (nx51070), .A0 (ram_223__6), .A1 (nx65538), .S0 (
             nx64214)) ;
    dffr reg_ram_222__6 (.Q (ram_222__6), .QB (\$dummy [1583]), .D (nx51080), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51081 (.Y (nx51080), .A0 (ram_222__6), .A1 (nx65538), .S0 (
             nx64218)) ;
    oai21 ix61288 (.Y (nx61287), .A0 (nx20026), .A1 (nx19948), .B0 (nx65108)) ;
    nand04 ix20027 (.Y (nx20026), .A0 (nx61290), .A1 (nx61298), .A2 (nx61306), .A3 (
           nx61314)) ;
    aoi22 ix61291 (.Y (nx61290), .A0 (ram_192__6), .A1 (nx64516), .B0 (
          ram_193__6), .B1 (nx64554)) ;
    dffr reg_ram_192__6 (.Q (ram_192__6), .QB (\$dummy [1584]), .D (nx51060), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51061 (.Y (nx51060), .A0 (ram_192__6), .A1 (nx65538), .S0 (
             nx64204)) ;
    dffr reg_ram_193__6 (.Q (ram_193__6), .QB (\$dummy [1585]), .D (nx51050), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51051 (.Y (nx51050), .A0 (ram_193__6), .A1 (nx65540), .S0 (
             nx64200)) ;
    aoi22 ix61299 (.Y (nx61298), .A0 (ram_195__6), .A1 (nx64592), .B0 (
          ram_194__6), .B1 (nx64630)) ;
    dffr reg_ram_195__6 (.Q (ram_195__6), .QB (\$dummy [1586]), .D (nx51030), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51031 (.Y (nx51030), .A0 (ram_195__6), .A1 (nx65540), .S0 (
             nx64192)) ;
    dffr reg_ram_194__6 (.Q (ram_194__6), .QB (\$dummy [1587]), .D (nx51040), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51041 (.Y (nx51040), .A0 (ram_194__6), .A1 (nx65540), .S0 (
             nx64196)) ;
    aoi22 ix61307 (.Y (nx61306), .A0 (ram_196__6), .A1 (nx64668), .B0 (
          ram_197__6), .B1 (nx64706)) ;
    dffr reg_ram_196__6 (.Q (ram_196__6), .QB (\$dummy [1588]), .D (nx51020), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51021 (.Y (nx51020), .A0 (ram_196__6), .A1 (nx65540), .S0 (
             nx64188)) ;
    dffr reg_ram_197__6 (.Q (ram_197__6), .QB (\$dummy [1589]), .D (nx51010), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51011 (.Y (nx51010), .A0 (ram_197__6), .A1 (nx65540), .S0 (
             nx64184)) ;
    aoi22 ix61315 (.Y (nx61314), .A0 (ram_199__6), .A1 (nx64744), .B0 (
          ram_198__6), .B1 (nx64782)) ;
    dffr reg_ram_199__6 (.Q (ram_199__6), .QB (\$dummy [1590]), .D (nx50990), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50991 (.Y (nx50990), .A0 (ram_199__6), .A1 (nx65540), .S0 (
             nx64176)) ;
    dffr reg_ram_198__6 (.Q (ram_198__6), .QB (\$dummy [1591]), .D (nx51000), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51001 (.Y (nx51000), .A0 (ram_198__6), .A1 (nx65540), .S0 (
             nx64180)) ;
    nand04 ix19949 (.Y (nx19948), .A0 (nx61323), .A1 (nx61331), .A2 (nx61339), .A3 (
           nx61347)) ;
    aoi22 ix61324 (.Y (nx61323), .A0 (ram_200__6), .A1 (nx64820), .B0 (
          ram_201__6), .B1 (nx64858)) ;
    dffr reg_ram_200__6 (.Q (ram_200__6), .QB (\$dummy [1592]), .D (nx50980), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50981 (.Y (nx50980), .A0 (ram_200__6), .A1 (nx65542), .S0 (
             nx64172)) ;
    dffr reg_ram_201__6 (.Q (ram_201__6), .QB (\$dummy [1593]), .D (nx50970), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50971 (.Y (nx50970), .A0 (ram_201__6), .A1 (nx65542), .S0 (
             nx64168)) ;
    aoi22 ix61332 (.Y (nx61331), .A0 (ram_203__6), .A1 (nx64896), .B0 (
          ram_202__6), .B1 (nx64934)) ;
    dffr reg_ram_203__6 (.Q (ram_203__6), .QB (\$dummy [1594]), .D (nx50950), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50951 (.Y (nx50950), .A0 (ram_203__6), .A1 (nx65542), .S0 (
             nx64160)) ;
    dffr reg_ram_202__6 (.Q (ram_202__6), .QB (\$dummy [1595]), .D (nx50960), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50961 (.Y (nx50960), .A0 (ram_202__6), .A1 (nx65542), .S0 (
             nx64164)) ;
    aoi22 ix61340 (.Y (nx61339), .A0 (ram_204__6), .A1 (nx64972), .B0 (
          ram_205__6), .B1 (nx65010)) ;
    dffr reg_ram_204__6 (.Q (ram_204__6), .QB (\$dummy [1596]), .D (nx50940), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50941 (.Y (nx50940), .A0 (ram_204__6), .A1 (nx65542), .S0 (
             nx64156)) ;
    dffr reg_ram_205__6 (.Q (ram_205__6), .QB (\$dummy [1597]), .D (nx50930), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50931 (.Y (nx50930), .A0 (ram_205__6), .A1 (nx65542), .S0 (
             nx64152)) ;
    aoi22 ix61348 (.Y (nx61347), .A0 (ram_207__6), .A1 (nx65048), .B0 (
          ram_206__6), .B1 (nx65086)) ;
    dffr reg_ram_207__6 (.Q (ram_207__6), .QB (\$dummy [1598]), .D (nx50910), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50911 (.Y (nx50910), .A0 (ram_207__6), .A1 (nx65542), .S0 (
             nx64144)) ;
    dffr reg_ram_206__6 (.Q (ram_206__6), .QB (\$dummy [1599]), .D (nx50920), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50921 (.Y (nx50920), .A0 (ram_206__6), .A1 (nx65544), .S0 (
             nx64148)) ;
    nand04 ix19871 (.Y (nx19870), .A0 (nx61356), .A1 (nx61424), .A2 (nx61492), .A3 (
           nx61560)) ;
    oai21 ix61357 (.Y (nx61356), .A0 (nx19860), .A1 (nx19782), .B0 (nx65112)) ;
    nand04 ix19861 (.Y (nx19860), .A0 (nx61359), .A1 (nx61367), .A2 (nx61375), .A3 (
           nx61383)) ;
    aoi22 ix61360 (.Y (nx61359), .A0 (ram_80__6), .A1 (nx64516), .B0 (ram_81__6)
          , .B1 (nx64554)) ;
    dffr reg_ram_80__6 (.Q (ram_80__6), .QB (\$dummy [1600]), .D (nx50900), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50901 (.Y (nx50900), .A0 (ram_80__6), .A1 (nx65544), .S0 (nx64134
             )) ;
    dffr reg_ram_81__6 (.Q (ram_81__6), .QB (\$dummy [1601]), .D (nx50890), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50891 (.Y (nx50890), .A0 (ram_81__6), .A1 (nx65544), .S0 (nx64130
             )) ;
    aoi22 ix61368 (.Y (nx61367), .A0 (ram_83__6), .A1 (nx64592), .B0 (ram_82__6)
          , .B1 (nx64630)) ;
    dffr reg_ram_83__6 (.Q (ram_83__6), .QB (\$dummy [1602]), .D (nx50870), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50871 (.Y (nx50870), .A0 (ram_83__6), .A1 (nx65544), .S0 (nx64122
             )) ;
    dffr reg_ram_82__6 (.Q (ram_82__6), .QB (\$dummy [1603]), .D (nx50880), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50881 (.Y (nx50880), .A0 (ram_82__6), .A1 (nx65544), .S0 (nx64126
             )) ;
    aoi22 ix61376 (.Y (nx61375), .A0 (ram_84__6), .A1 (nx64668), .B0 (ram_85__6)
          , .B1 (nx64706)) ;
    dffr reg_ram_84__6 (.Q (ram_84__6), .QB (\$dummy [1604]), .D (nx50860), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50861 (.Y (nx50860), .A0 (ram_84__6), .A1 (nx65544), .S0 (nx64118
             )) ;
    dffr reg_ram_85__6 (.Q (ram_85__6), .QB (\$dummy [1605]), .D (nx50850), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50851 (.Y (nx50850), .A0 (ram_85__6), .A1 (nx65544), .S0 (nx64114
             )) ;
    aoi22 ix61384 (.Y (nx61383), .A0 (ram_87__6), .A1 (nx64744), .B0 (ram_86__6)
          , .B1 (nx64782)) ;
    dffr reg_ram_87__6 (.Q (ram_87__6), .QB (\$dummy [1606]), .D (nx50830), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50831 (.Y (nx50830), .A0 (ram_87__6), .A1 (nx65546), .S0 (nx64106
             )) ;
    dffr reg_ram_86__6 (.Q (ram_86__6), .QB (\$dummy [1607]), .D (nx50840), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50841 (.Y (nx50840), .A0 (ram_86__6), .A1 (nx65546), .S0 (nx64110
             )) ;
    nand04 ix19783 (.Y (nx19782), .A0 (nx61392), .A1 (nx61400), .A2 (nx61408), .A3 (
           nx61416)) ;
    aoi22 ix61393 (.Y (nx61392), .A0 (ram_88__6), .A1 (nx64820), .B0 (ram_89__6)
          , .B1 (nx64858)) ;
    dffr reg_ram_88__6 (.Q (ram_88__6), .QB (\$dummy [1608]), .D (nx50820), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50821 (.Y (nx50820), .A0 (ram_88__6), .A1 (nx65546), .S0 (nx64102
             )) ;
    dffr reg_ram_89__6 (.Q (ram_89__6), .QB (\$dummy [1609]), .D (nx50810), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50811 (.Y (nx50810), .A0 (ram_89__6), .A1 (nx65546), .S0 (nx64098
             )) ;
    aoi22 ix61401 (.Y (nx61400), .A0 (ram_91__6), .A1 (nx64896), .B0 (ram_90__6)
          , .B1 (nx64934)) ;
    dffr reg_ram_91__6 (.Q (ram_91__6), .QB (\$dummy [1610]), .D (nx50790), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50791 (.Y (nx50790), .A0 (ram_91__6), .A1 (nx65546), .S0 (nx64090
             )) ;
    dffr reg_ram_90__6 (.Q (ram_90__6), .QB (\$dummy [1611]), .D (nx50800), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50801 (.Y (nx50800), .A0 (ram_90__6), .A1 (nx65546), .S0 (nx64094
             )) ;
    aoi22 ix61409 (.Y (nx61408), .A0 (ram_92__6), .A1 (nx64972), .B0 (ram_93__6)
          , .B1 (nx65010)) ;
    dffr reg_ram_92__6 (.Q (ram_92__6), .QB (\$dummy [1612]), .D (nx50780), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50781 (.Y (nx50780), .A0 (ram_92__6), .A1 (nx65546), .S0 (nx64086
             )) ;
    dffr reg_ram_93__6 (.Q (ram_93__6), .QB (\$dummy [1613]), .D (nx50770), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50771 (.Y (nx50770), .A0 (ram_93__6), .A1 (nx65548), .S0 (nx64082
             )) ;
    aoi22 ix61417 (.Y (nx61416), .A0 (ram_95__6), .A1 (nx65048), .B0 (ram_94__6)
          , .B1 (nx65086)) ;
    dffr reg_ram_95__6 (.Q (ram_95__6), .QB (\$dummy [1614]), .D (nx50750), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50751 (.Y (nx50750), .A0 (ram_95__6), .A1 (nx65548), .S0 (nx64074
             )) ;
    dffr reg_ram_94__6 (.Q (ram_94__6), .QB (\$dummy [1615]), .D (nx50760), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50761 (.Y (nx50760), .A0 (ram_94__6), .A1 (nx65548), .S0 (nx64078
             )) ;
    oai21 ix61425 (.Y (nx61424), .A0 (nx19698), .A1 (nx19620), .B0 (nx65116)) ;
    nand04 ix19699 (.Y (nx19698), .A0 (nx61427), .A1 (nx61435), .A2 (nx61443), .A3 (
           nx61451)) ;
    aoi22 ix61428 (.Y (nx61427), .A0 (ram_64__6), .A1 (nx64516), .B0 (ram_65__6)
          , .B1 (nx64554)) ;
    dffr reg_ram_64__6 (.Q (ram_64__6), .QB (\$dummy [1616]), .D (nx50740), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50741 (.Y (nx50740), .A0 (ram_64__6), .A1 (nx65548), .S0 (nx64064
             )) ;
    dffr reg_ram_65__6 (.Q (ram_65__6), .QB (\$dummy [1617]), .D (nx50730), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50731 (.Y (nx50730), .A0 (ram_65__6), .A1 (nx65548), .S0 (nx64060
             )) ;
    aoi22 ix61436 (.Y (nx61435), .A0 (ram_67__6), .A1 (nx64592), .B0 (ram_66__6)
          , .B1 (nx64630)) ;
    dffr reg_ram_67__6 (.Q (ram_67__6), .QB (\$dummy [1618]), .D (nx50710), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50711 (.Y (nx50710), .A0 (ram_67__6), .A1 (nx65548), .S0 (nx64052
             )) ;
    dffr reg_ram_66__6 (.Q (ram_66__6), .QB (\$dummy [1619]), .D (nx50720), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50721 (.Y (nx50720), .A0 (ram_66__6), .A1 (nx65548), .S0 (nx64056
             )) ;
    aoi22 ix61444 (.Y (nx61443), .A0 (ram_68__6), .A1 (nx64668), .B0 (ram_69__6)
          , .B1 (nx64706)) ;
    dffr reg_ram_68__6 (.Q (ram_68__6), .QB (\$dummy [1620]), .D (nx50700), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50701 (.Y (nx50700), .A0 (ram_68__6), .A1 (nx65550), .S0 (nx64048
             )) ;
    dffr reg_ram_69__6 (.Q (ram_69__6), .QB (\$dummy [1621]), .D (nx50690), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50691 (.Y (nx50690), .A0 (ram_69__6), .A1 (nx65550), .S0 (nx64044
             )) ;
    aoi22 ix61452 (.Y (nx61451), .A0 (ram_71__6), .A1 (nx64744), .B0 (ram_70__6)
          , .B1 (nx64782)) ;
    dffr reg_ram_71__6 (.Q (ram_71__6), .QB (\$dummy [1622]), .D (nx50670), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50671 (.Y (nx50670), .A0 (ram_71__6), .A1 (nx65550), .S0 (nx64036
             )) ;
    dffr reg_ram_70__6 (.Q (ram_70__6), .QB (\$dummy [1623]), .D (nx50680), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50681 (.Y (nx50680), .A0 (ram_70__6), .A1 (nx65550), .S0 (nx64040
             )) ;
    nand04 ix19621 (.Y (nx19620), .A0 (nx61460), .A1 (nx61468), .A2 (nx61476), .A3 (
           nx61484)) ;
    aoi22 ix61461 (.Y (nx61460), .A0 (ram_72__6), .A1 (nx64820), .B0 (ram_73__6)
          , .B1 (nx64858)) ;
    dffr reg_ram_72__6 (.Q (ram_72__6), .QB (\$dummy [1624]), .D (nx50660), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50661 (.Y (nx50660), .A0 (ram_72__6), .A1 (nx65550), .S0 (nx64032
             )) ;
    dffr reg_ram_73__6 (.Q (ram_73__6), .QB (\$dummy [1625]), .D (nx50650), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50651 (.Y (nx50650), .A0 (ram_73__6), .A1 (nx65550), .S0 (nx64028
             )) ;
    aoi22 ix61469 (.Y (nx61468), .A0 (ram_75__6), .A1 (nx64896), .B0 (ram_74__6)
          , .B1 (nx64934)) ;
    dffr reg_ram_75__6 (.Q (ram_75__6), .QB (\$dummy [1626]), .D (nx50630), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50631 (.Y (nx50630), .A0 (ram_75__6), .A1 (nx65550), .S0 (nx64020
             )) ;
    dffr reg_ram_74__6 (.Q (ram_74__6), .QB (\$dummy [1627]), .D (nx50640), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50641 (.Y (nx50640), .A0 (ram_74__6), .A1 (nx65552), .S0 (nx64024
             )) ;
    aoi22 ix61477 (.Y (nx61476), .A0 (ram_76__6), .A1 (nx64972), .B0 (ram_77__6)
          , .B1 (nx65010)) ;
    dffr reg_ram_76__6 (.Q (ram_76__6), .QB (\$dummy [1628]), .D (nx50620), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50621 (.Y (nx50620), .A0 (ram_76__6), .A1 (nx65552), .S0 (nx64016
             )) ;
    dffr reg_ram_77__6 (.Q (ram_77__6), .QB (\$dummy [1629]), .D (nx50610), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50611 (.Y (nx50610), .A0 (ram_77__6), .A1 (nx65552), .S0 (nx64012
             )) ;
    aoi22 ix61485 (.Y (nx61484), .A0 (ram_79__6), .A1 (nx65048), .B0 (ram_78__6)
          , .B1 (nx65086)) ;
    dffr reg_ram_79__6 (.Q (ram_79__6), .QB (\$dummy [1630]), .D (nx50590), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50591 (.Y (nx50590), .A0 (ram_79__6), .A1 (nx65552), .S0 (nx64004
             )) ;
    dffr reg_ram_78__6 (.Q (ram_78__6), .QB (\$dummy [1631]), .D (nx50600), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50601 (.Y (nx50600), .A0 (ram_78__6), .A1 (nx65552), .S0 (nx64008
             )) ;
    oai21 ix61493 (.Y (nx61492), .A0 (nx19534), .A1 (nx19456), .B0 (nx65120)) ;
    nand04 ix19535 (.Y (nx19534), .A0 (nx61495), .A1 (nx61503), .A2 (nx61511), .A3 (
           nx61519)) ;
    aoi22 ix61496 (.Y (nx61495), .A0 (ram_48__6), .A1 (nx64516), .B0 (ram_49__6)
          , .B1 (nx64554)) ;
    dffr reg_ram_48__6 (.Q (ram_48__6), .QB (\$dummy [1632]), .D (nx50580), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50581 (.Y (nx50580), .A0 (ram_48__6), .A1 (nx65552), .S0 (nx63994
             )) ;
    dffr reg_ram_49__6 (.Q (ram_49__6), .QB (\$dummy [1633]), .D (nx50570), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50571 (.Y (nx50570), .A0 (ram_49__6), .A1 (nx65552), .S0 (nx63990
             )) ;
    aoi22 ix61504 (.Y (nx61503), .A0 (ram_51__6), .A1 (nx64592), .B0 (ram_50__6)
          , .B1 (nx64630)) ;
    dffr reg_ram_51__6 (.Q (ram_51__6), .QB (\$dummy [1634]), .D (nx50550), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50551 (.Y (nx50550), .A0 (ram_51__6), .A1 (nx65554), .S0 (nx63982
             )) ;
    dffr reg_ram_50__6 (.Q (ram_50__6), .QB (\$dummy [1635]), .D (nx50560), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50561 (.Y (nx50560), .A0 (ram_50__6), .A1 (nx65554), .S0 (nx63986
             )) ;
    aoi22 ix61512 (.Y (nx61511), .A0 (ram_52__6), .A1 (nx64668), .B0 (ram_53__6)
          , .B1 (nx64706)) ;
    dffr reg_ram_52__6 (.Q (ram_52__6), .QB (\$dummy [1636]), .D (nx50540), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50541 (.Y (nx50540), .A0 (ram_52__6), .A1 (nx65554), .S0 (nx63978
             )) ;
    dffr reg_ram_53__6 (.Q (ram_53__6), .QB (\$dummy [1637]), .D (nx50530), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50531 (.Y (nx50530), .A0 (ram_53__6), .A1 (nx65554), .S0 (nx63974
             )) ;
    aoi22 ix61520 (.Y (nx61519), .A0 (ram_55__6), .A1 (nx64744), .B0 (ram_54__6)
          , .B1 (nx64782)) ;
    dffr reg_ram_55__6 (.Q (ram_55__6), .QB (\$dummy [1638]), .D (nx50510), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50511 (.Y (nx50510), .A0 (ram_55__6), .A1 (nx65554), .S0 (nx63966
             )) ;
    dffr reg_ram_54__6 (.Q (ram_54__6), .QB (\$dummy [1639]), .D (nx50520), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50521 (.Y (nx50520), .A0 (ram_54__6), .A1 (nx65554), .S0 (nx63970
             )) ;
    nand04 ix19457 (.Y (nx19456), .A0 (nx61528), .A1 (nx61536), .A2 (nx61544), .A3 (
           nx61552)) ;
    aoi22 ix61529 (.Y (nx61528), .A0 (ram_56__6), .A1 (nx64820), .B0 (ram_57__6)
          , .B1 (nx64858)) ;
    dffr reg_ram_56__6 (.Q (ram_56__6), .QB (\$dummy [1640]), .D (nx50500), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50501 (.Y (nx50500), .A0 (ram_56__6), .A1 (nx65554), .S0 (nx63962
             )) ;
    dffr reg_ram_57__6 (.Q (ram_57__6), .QB (\$dummy [1641]), .D (nx50490), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50491 (.Y (nx50490), .A0 (ram_57__6), .A1 (nx65556), .S0 (nx63958
             )) ;
    aoi22 ix61537 (.Y (nx61536), .A0 (ram_59__6), .A1 (nx64896), .B0 (ram_58__6)
          , .B1 (nx64934)) ;
    dffr reg_ram_59__6 (.Q (ram_59__6), .QB (\$dummy [1642]), .D (nx50470), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50471 (.Y (nx50470), .A0 (ram_59__6), .A1 (nx65556), .S0 (nx63950
             )) ;
    dffr reg_ram_58__6 (.Q (ram_58__6), .QB (\$dummy [1643]), .D (nx50480), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50481 (.Y (nx50480), .A0 (ram_58__6), .A1 (nx65556), .S0 (nx63954
             )) ;
    aoi22 ix61545 (.Y (nx61544), .A0 (ram_60__6), .A1 (nx64972), .B0 (ram_61__6)
          , .B1 (nx65010)) ;
    dffr reg_ram_60__6 (.Q (ram_60__6), .QB (\$dummy [1644]), .D (nx50460), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50461 (.Y (nx50460), .A0 (ram_60__6), .A1 (nx65556), .S0 (nx63946
             )) ;
    dffr reg_ram_61__6 (.Q (ram_61__6), .QB (\$dummy [1645]), .D (nx50450), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50451 (.Y (nx50450), .A0 (ram_61__6), .A1 (nx65556), .S0 (nx63942
             )) ;
    aoi22 ix61553 (.Y (nx61552), .A0 (ram_63__6), .A1 (nx65048), .B0 (ram_62__6)
          , .B1 (nx65086)) ;
    dffr reg_ram_63__6 (.Q (ram_63__6), .QB (\$dummy [1646]), .D (nx50430), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50431 (.Y (nx50430), .A0 (ram_63__6), .A1 (nx65556), .S0 (nx63934
             )) ;
    dffr reg_ram_62__6 (.Q (ram_62__6), .QB (\$dummy [1647]), .D (nx50440), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50441 (.Y (nx50440), .A0 (ram_62__6), .A1 (nx65556), .S0 (nx63938
             )) ;
    oai21 ix61561 (.Y (nx61560), .A0 (nx19372), .A1 (nx19294), .B0 (nx65124)) ;
    nand04 ix19373 (.Y (nx19372), .A0 (nx61563), .A1 (nx61571), .A2 (nx61579), .A3 (
           nx61587)) ;
    aoi22 ix61564 (.Y (nx61563), .A0 (ram_32__6), .A1 (nx64516), .B0 (ram_33__6)
          , .B1 (nx64554)) ;
    dffr reg_ram_32__6 (.Q (ram_32__6), .QB (\$dummy [1648]), .D (nx50420), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50421 (.Y (nx50420), .A0 (ram_32__6), .A1 (nx65558), .S0 (nx63924
             )) ;
    dffr reg_ram_33__6 (.Q (ram_33__6), .QB (\$dummy [1649]), .D (nx50410), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50411 (.Y (nx50410), .A0 (ram_33__6), .A1 (nx65558), .S0 (nx63920
             )) ;
    aoi22 ix61572 (.Y (nx61571), .A0 (ram_35__6), .A1 (nx64592), .B0 (ram_34__6)
          , .B1 (nx64630)) ;
    dffr reg_ram_35__6 (.Q (ram_35__6), .QB (\$dummy [1650]), .D (nx50390), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50391 (.Y (nx50390), .A0 (ram_35__6), .A1 (nx65558), .S0 (nx63912
             )) ;
    dffr reg_ram_34__6 (.Q (ram_34__6), .QB (\$dummy [1651]), .D (nx50400), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50401 (.Y (nx50400), .A0 (ram_34__6), .A1 (nx65558), .S0 (nx63916
             )) ;
    aoi22 ix61580 (.Y (nx61579), .A0 (ram_36__6), .A1 (nx64668), .B0 (ram_37__6)
          , .B1 (nx64706)) ;
    dffr reg_ram_36__6 (.Q (ram_36__6), .QB (\$dummy [1652]), .D (nx50380), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50381 (.Y (nx50380), .A0 (ram_36__6), .A1 (nx65558), .S0 (nx63908
             )) ;
    dffr reg_ram_37__6 (.Q (ram_37__6), .QB (\$dummy [1653]), .D (nx50370), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50371 (.Y (nx50370), .A0 (ram_37__6), .A1 (nx65558), .S0 (nx63904
             )) ;
    aoi22 ix61588 (.Y (nx61587), .A0 (ram_39__6), .A1 (nx64744), .B0 (ram_38__6)
          , .B1 (nx64782)) ;
    dffr reg_ram_39__6 (.Q (ram_39__6), .QB (\$dummy [1654]), .D (nx50350), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50351 (.Y (nx50350), .A0 (ram_39__6), .A1 (nx65558), .S0 (nx63896
             )) ;
    dffr reg_ram_38__6 (.Q (ram_38__6), .QB (\$dummy [1655]), .D (nx50360), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50361 (.Y (nx50360), .A0 (ram_38__6), .A1 (nx65560), .S0 (nx63900
             )) ;
    nand04 ix19295 (.Y (nx19294), .A0 (nx61596), .A1 (nx61604), .A2 (nx61612), .A3 (
           nx61620)) ;
    aoi22 ix61597 (.Y (nx61596), .A0 (ram_40__6), .A1 (nx64820), .B0 (ram_41__6)
          , .B1 (nx64858)) ;
    dffr reg_ram_40__6 (.Q (ram_40__6), .QB (\$dummy [1656]), .D (nx50340), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50341 (.Y (nx50340), .A0 (ram_40__6), .A1 (nx65560), .S0 (nx63892
             )) ;
    dffr reg_ram_41__6 (.Q (ram_41__6), .QB (\$dummy [1657]), .D (nx50330), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50331 (.Y (nx50330), .A0 (ram_41__6), .A1 (nx65560), .S0 (nx63888
             )) ;
    aoi22 ix61605 (.Y (nx61604), .A0 (ram_43__6), .A1 (nx64896), .B0 (ram_42__6)
          , .B1 (nx64934)) ;
    dffr reg_ram_43__6 (.Q (ram_43__6), .QB (\$dummy [1658]), .D (nx50310), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50311 (.Y (nx50310), .A0 (ram_43__6), .A1 (nx65560), .S0 (nx63880
             )) ;
    dffr reg_ram_42__6 (.Q (ram_42__6), .QB (\$dummy [1659]), .D (nx50320), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50321 (.Y (nx50320), .A0 (ram_42__6), .A1 (nx65560), .S0 (nx63884
             )) ;
    aoi22 ix61613 (.Y (nx61612), .A0 (ram_44__6), .A1 (nx64972), .B0 (ram_45__6)
          , .B1 (nx65010)) ;
    dffr reg_ram_44__6 (.Q (ram_44__6), .QB (\$dummy [1660]), .D (nx50300), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50301 (.Y (nx50300), .A0 (ram_44__6), .A1 (nx65560), .S0 (nx63876
             )) ;
    dffr reg_ram_45__6 (.Q (ram_45__6), .QB (\$dummy [1661]), .D (nx50290), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50291 (.Y (nx50290), .A0 (ram_45__6), .A1 (nx65560), .S0 (nx63872
             )) ;
    aoi22 ix61621 (.Y (nx61620), .A0 (ram_47__6), .A1 (nx65048), .B0 (ram_46__6)
          , .B1 (nx65086)) ;
    dffr reg_ram_47__6 (.Q (ram_47__6), .QB (\$dummy [1662]), .D (nx50270), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50271 (.Y (nx50270), .A0 (ram_47__6), .A1 (nx65562), .S0 (nx63864
             )) ;
    dffr reg_ram_46__6 (.Q (ram_46__6), .QB (\$dummy [1663]), .D (nx50280), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50281 (.Y (nx50280), .A0 (ram_46__6), .A1 (nx65562), .S0 (nx63868
             )) ;
    nand04 ix19215 (.Y (nx19214), .A0 (nx61629), .A1 (nx61697), .A2 (nx61765), .A3 (
           nx61833)) ;
    oai21 ix61630 (.Y (nx61629), .A0 (nx19204), .A1 (nx19126), .B0 (nx65128)) ;
    nand04 ix19205 (.Y (nx19204), .A0 (nx61632), .A1 (nx61640), .A2 (nx61648), .A3 (
           nx61656)) ;
    aoi22 ix61633 (.Y (nx61632), .A0 (ram_16__6), .A1 (nx64518), .B0 (ram_17__6)
          , .B1 (nx64556)) ;
    dffr reg_ram_16__6 (.Q (ram_16__6), .QB (\$dummy [1664]), .D (nx50260), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50261 (.Y (nx50260), .A0 (ram_16__6), .A1 (nx65562), .S0 (nx63854
             )) ;
    dffr reg_ram_17__6 (.Q (ram_17__6), .QB (\$dummy [1665]), .D (nx50250), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50251 (.Y (nx50250), .A0 (ram_17__6), .A1 (nx65562), .S0 (nx63850
             )) ;
    aoi22 ix61641 (.Y (nx61640), .A0 (ram_19__6), .A1 (nx64594), .B0 (ram_18__6)
          , .B1 (nx64632)) ;
    dffr reg_ram_19__6 (.Q (ram_19__6), .QB (\$dummy [1666]), .D (nx50230), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50231 (.Y (nx50230), .A0 (ram_19__6), .A1 (nx65562), .S0 (nx63842
             )) ;
    dffr reg_ram_18__6 (.Q (ram_18__6), .QB (\$dummy [1667]), .D (nx50240), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50241 (.Y (nx50240), .A0 (ram_18__6), .A1 (nx65562), .S0 (nx63846
             )) ;
    aoi22 ix61649 (.Y (nx61648), .A0 (ram_20__6), .A1 (nx64670), .B0 (ram_21__6)
          , .B1 (nx64708)) ;
    dffr reg_ram_20__6 (.Q (ram_20__6), .QB (\$dummy [1668]), .D (nx50220), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50221 (.Y (nx50220), .A0 (ram_20__6), .A1 (nx65562), .S0 (nx63838
             )) ;
    dffr reg_ram_21__6 (.Q (ram_21__6), .QB (\$dummy [1669]), .D (nx50210), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50211 (.Y (nx50210), .A0 (ram_21__6), .A1 (nx65564), .S0 (nx63834
             )) ;
    aoi22 ix61657 (.Y (nx61656), .A0 (ram_23__6), .A1 (nx64746), .B0 (ram_22__6)
          , .B1 (nx64784)) ;
    dffr reg_ram_23__6 (.Q (ram_23__6), .QB (\$dummy [1670]), .D (nx50190), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50191 (.Y (nx50190), .A0 (ram_23__6), .A1 (nx65564), .S0 (nx63826
             )) ;
    dffr reg_ram_22__6 (.Q (ram_22__6), .QB (\$dummy [1671]), .D (nx50200), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50201 (.Y (nx50200), .A0 (ram_22__6), .A1 (nx65564), .S0 (nx63830
             )) ;
    nand04 ix19127 (.Y (nx19126), .A0 (nx61665), .A1 (nx61673), .A2 (nx61681), .A3 (
           nx61689)) ;
    aoi22 ix61666 (.Y (nx61665), .A0 (ram_24__6), .A1 (nx64822), .B0 (ram_25__6)
          , .B1 (nx64860)) ;
    dffr reg_ram_24__6 (.Q (ram_24__6), .QB (\$dummy [1672]), .D (nx50180), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50181 (.Y (nx50180), .A0 (ram_24__6), .A1 (nx65564), .S0 (nx63822
             )) ;
    dffr reg_ram_25__6 (.Q (ram_25__6), .QB (\$dummy [1673]), .D (nx50170), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50171 (.Y (nx50170), .A0 (ram_25__6), .A1 (nx65564), .S0 (nx63818
             )) ;
    aoi22 ix61674 (.Y (nx61673), .A0 (ram_27__6), .A1 (nx64898), .B0 (ram_26__6)
          , .B1 (nx64936)) ;
    dffr reg_ram_27__6 (.Q (ram_27__6), .QB (\$dummy [1674]), .D (nx50150), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50151 (.Y (nx50150), .A0 (ram_27__6), .A1 (nx65564), .S0 (nx63810
             )) ;
    dffr reg_ram_26__6 (.Q (ram_26__6), .QB (\$dummy [1675]), .D (nx50160), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50161 (.Y (nx50160), .A0 (ram_26__6), .A1 (nx65564), .S0 (nx63814
             )) ;
    aoi22 ix61682 (.Y (nx61681), .A0 (ram_28__6), .A1 (nx64974), .B0 (ram_29__6)
          , .B1 (nx65012)) ;
    dffr reg_ram_28__6 (.Q (ram_28__6), .QB (\$dummy [1676]), .D (nx50140), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50141 (.Y (nx50140), .A0 (ram_28__6), .A1 (nx65566), .S0 (nx63806
             )) ;
    dffr reg_ram_29__6 (.Q (ram_29__6), .QB (\$dummy [1677]), .D (nx50130), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50131 (.Y (nx50130), .A0 (ram_29__6), .A1 (nx65566), .S0 (nx63802
             )) ;
    aoi22 ix61690 (.Y (nx61689), .A0 (ram_31__6), .A1 (nx65050), .B0 (ram_30__6)
          , .B1 (nx65088)) ;
    dffr reg_ram_31__6 (.Q (ram_31__6), .QB (\$dummy [1678]), .D (nx50110), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50111 (.Y (nx50110), .A0 (ram_31__6), .A1 (nx65566), .S0 (nx63794
             )) ;
    dffr reg_ram_30__6 (.Q (ram_30__6), .QB (\$dummy [1679]), .D (nx50120), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50121 (.Y (nx50120), .A0 (ram_30__6), .A1 (nx65566), .S0 (nx63798
             )) ;
    oai21 ix61698 (.Y (nx61697), .A0 (nx19042), .A1 (nx18964), .B0 (nx65144)) ;
    nand04 ix19043 (.Y (nx19042), .A0 (nx61700), .A1 (nx61708), .A2 (nx61716), .A3 (
           nx61724)) ;
    aoi22 ix61701 (.Y (nx61700), .A0 (ram_0__6), .A1 (nx64518), .B0 (ram_1__6), 
          .B1 (nx64556)) ;
    dffr reg_ram_0__6 (.Q (ram_0__6), .QB (\$dummy [1680]), .D (nx50100), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50101 (.Y (nx50100), .A0 (nx65566), .A1 (ram_0__6), .S0 (nx65132)
             ) ;
    dffr reg_ram_1__6 (.Q (ram_1__6), .QB (\$dummy [1681]), .D (nx50090), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50091 (.Y (nx50090), .A0 (nx65566), .A1 (ram_1__6), .S0 (nx65146)
             ) ;
    aoi22 ix61709 (.Y (nx61708), .A0 (ram_3__6), .A1 (nx64594), .B0 (ram_2__6), 
          .B1 (nx64632)) ;
    dffr reg_ram_3__6 (.Q (ram_3__6), .QB (\$dummy [1682]), .D (nx50070), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50071 (.Y (nx50070), .A0 (nx65566), .A1 (ram_3__6), .S0 (nx65150)
             ) ;
    dffr reg_ram_2__6 (.Q (ram_2__6), .QB (\$dummy [1683]), .D (nx50080), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50081 (.Y (nx50080), .A0 (nx65568), .A1 (ram_2__6), .S0 (nx65154)
             ) ;
    aoi22 ix61717 (.Y (nx61716), .A0 (ram_4__6), .A1 (nx64670), .B0 (ram_5__6), 
          .B1 (nx64708)) ;
    dffr reg_ram_4__6 (.Q (ram_4__6), .QB (\$dummy [1684]), .D (nx50060), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50061 (.Y (nx50060), .A0 (nx65568), .A1 (ram_4__6), .S0 (nx65158)
             ) ;
    dffr reg_ram_5__6 (.Q (ram_5__6), .QB (\$dummy [1685]), .D (nx50050), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50051 (.Y (nx50050), .A0 (nx65568), .A1 (ram_5__6), .S0 (nx65162)
             ) ;
    aoi22 ix61725 (.Y (nx61724), .A0 (ram_7__6), .A1 (nx64746), .B0 (ram_6__6), 
          .B1 (nx64784)) ;
    dffr reg_ram_7__6 (.Q (ram_7__6), .QB (\$dummy [1686]), .D (nx50030), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50031 (.Y (nx50030), .A0 (nx65568), .A1 (ram_7__6), .S0 (nx65166)
             ) ;
    dffr reg_ram_6__6 (.Q (ram_6__6), .QB (\$dummy [1687]), .D (nx50040), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50041 (.Y (nx50040), .A0 (nx65568), .A1 (ram_6__6), .S0 (nx65170)
             ) ;
    nand04 ix18965 (.Y (nx18964), .A0 (nx61733), .A1 (nx61741), .A2 (nx61749), .A3 (
           nx61757)) ;
    aoi22 ix61734 (.Y (nx61733), .A0 (ram_8__6), .A1 (nx64822), .B0 (ram_9__6), 
          .B1 (nx64860)) ;
    dffr reg_ram_8__6 (.Q (ram_8__6), .QB (\$dummy [1688]), .D (nx50020), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50021 (.Y (nx50020), .A0 (nx65568), .A1 (ram_8__6), .S0 (nx65174)
             ) ;
    dffr reg_ram_9__6 (.Q (ram_9__6), .QB (\$dummy [1689]), .D (nx50010), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50011 (.Y (nx50010), .A0 (nx65568), .A1 (ram_9__6), .S0 (nx65178)
             ) ;
    aoi22 ix61742 (.Y (nx61741), .A0 (ram_11__6), .A1 (nx64898), .B0 (ram_10__6)
          , .B1 (nx64936)) ;
    dffr reg_ram_11__6 (.Q (ram_11__6), .QB (\$dummy [1690]), .D (nx49990), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49991 (.Y (nx49990), .A0 (nx65570), .A1 (ram_11__6), .S0 (nx65182
             )) ;
    dffr reg_ram_10__6 (.Q (ram_10__6), .QB (\$dummy [1691]), .D (nx50000), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix50001 (.Y (nx50000), .A0 (nx65570), .A1 (ram_10__6), .S0 (nx65186
             )) ;
    aoi22 ix61750 (.Y (nx61749), .A0 (ram_12__6), .A1 (nx64974), .B0 (ram_13__6)
          , .B1 (nx65012)) ;
    dffr reg_ram_12__6 (.Q (ram_12__6), .QB (\$dummy [1692]), .D (nx49980), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49981 (.Y (nx49980), .A0 (nx65570), .A1 (ram_12__6), .S0 (nx65190
             )) ;
    dffr reg_ram_13__6 (.Q (ram_13__6), .QB (\$dummy [1693]), .D (nx49970), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49971 (.Y (nx49970), .A0 (nx65570), .A1 (ram_13__6), .S0 (nx65194
             )) ;
    aoi22 ix61758 (.Y (nx61757), .A0 (ram_15__6), .A1 (nx65050), .B0 (ram_14__6)
          , .B1 (nx65088)) ;
    dffr reg_ram_15__6 (.Q (ram_15__6), .QB (\$dummy [1694]), .D (nx49950), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49951 (.Y (nx49950), .A0 (nx65570), .A1 (ram_15__6), .S0 (nx65198
             )) ;
    dffr reg_ram_14__6 (.Q (ram_14__6), .QB (\$dummy [1695]), .D (nx49960), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49961 (.Y (nx49960), .A0 (nx65570), .A1 (ram_14__6), .S0 (nx65202
             )) ;
    oai21 ix61766 (.Y (nx61765), .A0 (nx18878), .A1 (nx18800), .B0 (nx65206)) ;
    nand04 ix18879 (.Y (nx18878), .A0 (nx61768), .A1 (nx61776), .A2 (nx61784), .A3 (
           nx61792)) ;
    aoi22 ix61769 (.Y (nx61768), .A0 (ram_96__6), .A1 (nx64518), .B0 (ram_97__6)
          , .B1 (nx64556)) ;
    dffr reg_ram_96__6 (.Q (ram_96__6), .QB (\$dummy [1696]), .D (nx49940), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49941 (.Y (nx49940), .A0 (ram_96__6), .A1 (nx65570), .S0 (nx63784
             )) ;
    dffr reg_ram_97__6 (.Q (ram_97__6), .QB (\$dummy [1697]), .D (nx49930), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49931 (.Y (nx49930), .A0 (ram_97__6), .A1 (nx65572), .S0 (nx63780
             )) ;
    aoi22 ix61777 (.Y (nx61776), .A0 (ram_99__6), .A1 (nx64594), .B0 (ram_98__6)
          , .B1 (nx64632)) ;
    dffr reg_ram_99__6 (.Q (ram_99__6), .QB (\$dummy [1698]), .D (nx49910), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49911 (.Y (nx49910), .A0 (ram_99__6), .A1 (nx65572), .S0 (nx63772
             )) ;
    dffr reg_ram_98__6 (.Q (ram_98__6), .QB (\$dummy [1699]), .D (nx49920), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49921 (.Y (nx49920), .A0 (ram_98__6), .A1 (nx65572), .S0 (nx63776
             )) ;
    aoi22 ix61785 (.Y (nx61784), .A0 (ram_100__6), .A1 (nx64670), .B0 (
          ram_101__6), .B1 (nx64708)) ;
    dffr reg_ram_100__6 (.Q (ram_100__6), .QB (\$dummy [1700]), .D (nx49900), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49901 (.Y (nx49900), .A0 (ram_100__6), .A1 (nx65572), .S0 (
             nx63768)) ;
    dffr reg_ram_101__6 (.Q (ram_101__6), .QB (\$dummy [1701]), .D (nx49890), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49891 (.Y (nx49890), .A0 (ram_101__6), .A1 (nx65572), .S0 (
             nx63764)) ;
    aoi22 ix61793 (.Y (nx61792), .A0 (ram_103__6), .A1 (nx64746), .B0 (
          ram_102__6), .B1 (nx64784)) ;
    dffr reg_ram_103__6 (.Q (ram_103__6), .QB (\$dummy [1702]), .D (nx49870), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49871 (.Y (nx49870), .A0 (ram_103__6), .A1 (nx65572), .S0 (
             nx63756)) ;
    dffr reg_ram_102__6 (.Q (ram_102__6), .QB (\$dummy [1703]), .D (nx49880), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49881 (.Y (nx49880), .A0 (ram_102__6), .A1 (nx65572), .S0 (
             nx63760)) ;
    nand04 ix18801 (.Y (nx18800), .A0 (nx61801), .A1 (nx61809), .A2 (nx61817), .A3 (
           nx61825)) ;
    aoi22 ix61802 (.Y (nx61801), .A0 (ram_104__6), .A1 (nx64822), .B0 (
          ram_105__6), .B1 (nx64860)) ;
    dffr reg_ram_104__6 (.Q (ram_104__6), .QB (\$dummy [1704]), .D (nx49860), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49861 (.Y (nx49860), .A0 (ram_104__6), .A1 (nx65574), .S0 (
             nx63752)) ;
    dffr reg_ram_105__6 (.Q (ram_105__6), .QB (\$dummy [1705]), .D (nx49850), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49851 (.Y (nx49850), .A0 (ram_105__6), .A1 (nx65574), .S0 (
             nx63748)) ;
    aoi22 ix61810 (.Y (nx61809), .A0 (ram_107__6), .A1 (nx64898), .B0 (
          ram_106__6), .B1 (nx64936)) ;
    dffr reg_ram_107__6 (.Q (ram_107__6), .QB (\$dummy [1706]), .D (nx49830), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49831 (.Y (nx49830), .A0 (ram_107__6), .A1 (nx65574), .S0 (
             nx63740)) ;
    dffr reg_ram_106__6 (.Q (ram_106__6), .QB (\$dummy [1707]), .D (nx49840), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49841 (.Y (nx49840), .A0 (ram_106__6), .A1 (nx65574), .S0 (
             nx63744)) ;
    aoi22 ix61818 (.Y (nx61817), .A0 (ram_108__6), .A1 (nx64974), .B0 (
          ram_109__6), .B1 (nx65012)) ;
    dffr reg_ram_108__6 (.Q (ram_108__6), .QB (\$dummy [1708]), .D (nx49820), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49821 (.Y (nx49820), .A0 (ram_108__6), .A1 (nx65574), .S0 (
             nx63736)) ;
    dffr reg_ram_109__6 (.Q (ram_109__6), .QB (\$dummy [1709]), .D (nx49810), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49811 (.Y (nx49810), .A0 (ram_109__6), .A1 (nx65574), .S0 (
             nx63732)) ;
    aoi22 ix61826 (.Y (nx61825), .A0 (ram_111__6), .A1 (nx65050), .B0 (
          ram_110__6), .B1 (nx65088)) ;
    dffr reg_ram_111__6 (.Q (ram_111__6), .QB (\$dummy [1710]), .D (nx49790), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49791 (.Y (nx49790), .A0 (ram_111__6), .A1 (nx65574), .S0 (
             nx63724)) ;
    dffr reg_ram_110__6 (.Q (ram_110__6), .QB (\$dummy [1711]), .D (nx49800), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49801 (.Y (nx49800), .A0 (ram_110__6), .A1 (nx65576), .S0 (
             nx63728)) ;
    oai21 ix61834 (.Y (nx61833), .A0 (nx18716), .A1 (nx18638), .B0 (nx65210)) ;
    nand04 ix18717 (.Y (nx18716), .A0 (nx61836), .A1 (nx61844), .A2 (nx61852), .A3 (
           nx61860)) ;
    aoi22 ix61837 (.Y (nx61836), .A0 (ram_112__6), .A1 (nx64518), .B0 (
          ram_113__6), .B1 (nx64556)) ;
    dffr reg_ram_112__6 (.Q (ram_112__6), .QB (\$dummy [1712]), .D (nx49780), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49781 (.Y (nx49780), .A0 (ram_112__6), .A1 (nx65576), .S0 (
             nx63714)) ;
    dffr reg_ram_113__6 (.Q (ram_113__6), .QB (\$dummy [1713]), .D (nx49770), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49771 (.Y (nx49770), .A0 (ram_113__6), .A1 (nx65576), .S0 (
             nx63710)) ;
    aoi22 ix61845 (.Y (nx61844), .A0 (ram_115__6), .A1 (nx64594), .B0 (
          ram_114__6), .B1 (nx64632)) ;
    dffr reg_ram_115__6 (.Q (ram_115__6), .QB (\$dummy [1714]), .D (nx49750), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49751 (.Y (nx49750), .A0 (ram_115__6), .A1 (nx65576), .S0 (
             nx63702)) ;
    dffr reg_ram_114__6 (.Q (ram_114__6), .QB (\$dummy [1715]), .D (nx49760), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49761 (.Y (nx49760), .A0 (ram_114__6), .A1 (nx65576), .S0 (
             nx63706)) ;
    aoi22 ix61853 (.Y (nx61852), .A0 (ram_116__6), .A1 (nx64670), .B0 (
          ram_117__6), .B1 (nx64708)) ;
    dffr reg_ram_116__6 (.Q (ram_116__6), .QB (\$dummy [1716]), .D (nx49740), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49741 (.Y (nx49740), .A0 (ram_116__6), .A1 (nx65576), .S0 (
             nx63698)) ;
    dffr reg_ram_117__6 (.Q (ram_117__6), .QB (\$dummy [1717]), .D (nx49730), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49731 (.Y (nx49730), .A0 (ram_117__6), .A1 (nx65576), .S0 (
             nx63694)) ;
    aoi22 ix61861 (.Y (nx61860), .A0 (ram_119__6), .A1 (nx64746), .B0 (
          ram_118__6), .B1 (nx64784)) ;
    dffr reg_ram_119__6 (.Q (ram_119__6), .QB (\$dummy [1718]), .D (nx49710), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49711 (.Y (nx49710), .A0 (ram_119__6), .A1 (nx65578), .S0 (
             nx63686)) ;
    dffr reg_ram_118__6 (.Q (ram_118__6), .QB (\$dummy [1719]), .D (nx49720), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49721 (.Y (nx49720), .A0 (ram_118__6), .A1 (nx65578), .S0 (
             nx63690)) ;
    nand04 ix18639 (.Y (nx18638), .A0 (nx61869), .A1 (nx61877), .A2 (nx61885), .A3 (
           nx61893)) ;
    aoi22 ix61870 (.Y (nx61869), .A0 (ram_120__6), .A1 (nx64822), .B0 (
          ram_121__6), .B1 (nx64860)) ;
    dffr reg_ram_120__6 (.Q (ram_120__6), .QB (\$dummy [1720]), .D (nx49700), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49701 (.Y (nx49700), .A0 (ram_120__6), .A1 (nx65578), .S0 (
             nx63682)) ;
    dffr reg_ram_121__6 (.Q (ram_121__6), .QB (\$dummy [1721]), .D (nx49690), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49691 (.Y (nx49690), .A0 (ram_121__6), .A1 (nx65578), .S0 (
             nx63678)) ;
    aoi22 ix61878 (.Y (nx61877), .A0 (ram_123__6), .A1 (nx64898), .B0 (
          ram_122__6), .B1 (nx64936)) ;
    dffr reg_ram_123__6 (.Q (ram_123__6), .QB (\$dummy [1722]), .D (nx49670), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49671 (.Y (nx49670), .A0 (ram_123__6), .A1 (nx65578), .S0 (
             nx63670)) ;
    dffr reg_ram_122__6 (.Q (ram_122__6), .QB (\$dummy [1723]), .D (nx49680), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49681 (.Y (nx49680), .A0 (ram_122__6), .A1 (nx65578), .S0 (
             nx63674)) ;
    aoi22 ix61886 (.Y (nx61885), .A0 (ram_124__6), .A1 (nx64974), .B0 (
          ram_125__6), .B1 (nx65012)) ;
    dffr reg_ram_124__6 (.Q (ram_124__6), .QB (\$dummy [1724]), .D (nx49660), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49661 (.Y (nx49660), .A0 (ram_124__6), .A1 (nx65578), .S0 (
             nx63666)) ;
    dffr reg_ram_125__6 (.Q (ram_125__6), .QB (\$dummy [1725]), .D (nx49650), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49651 (.Y (nx49650), .A0 (ram_125__6), .A1 (nx65580), .S0 (
             nx63662)) ;
    aoi22 ix61894 (.Y (nx61893), .A0 (ram_127__6), .A1 (nx65050), .B0 (
          ram_126__6), .B1 (nx65088)) ;
    dffr reg_ram_127__6 (.Q (ram_127__6), .QB (\$dummy [1726]), .D (nx49630), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49631 (.Y (nx49630), .A0 (ram_127__6), .A1 (nx65580), .S0 (
             nx63654)) ;
    dffr reg_ram_126__6 (.Q (ram_126__6), .QB (\$dummy [1727]), .D (nx49640), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49641 (.Y (nx49640), .A0 (ram_126__6), .A1 (nx65580), .S0 (
             nx63658)) ;
    nand04 ix18561 (.Y (nx18560), .A0 (nx61902), .A1 (nx61970), .A2 (nx62038), .A3 (
           nx62106)) ;
    oai21 ix61903 (.Y (nx61902), .A0 (nx18550), .A1 (nx18472), .B0 (nx65214)) ;
    nand04 ix18551 (.Y (nx18550), .A0 (nx61905), .A1 (nx61913), .A2 (nx61921), .A3 (
           nx61929)) ;
    aoi22 ix61906 (.Y (nx61905), .A0 (ram_128__6), .A1 (nx64518), .B0 (
          ram_129__6), .B1 (nx64556)) ;
    dffr reg_ram_128__6 (.Q (ram_128__6), .QB (\$dummy [1728]), .D (nx49620), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49621 (.Y (nx49620), .A0 (ram_128__6), .A1 (nx65580), .S0 (
             nx63644)) ;
    dffr reg_ram_129__6 (.Q (ram_129__6), .QB (\$dummy [1729]), .D (nx49610), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49611 (.Y (nx49610), .A0 (ram_129__6), .A1 (nx65580), .S0 (
             nx63640)) ;
    aoi22 ix61914 (.Y (nx61913), .A0 (ram_131__6), .A1 (nx64594), .B0 (
          ram_130__6), .B1 (nx64632)) ;
    dffr reg_ram_131__6 (.Q (ram_131__6), .QB (\$dummy [1730]), .D (nx49590), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49591 (.Y (nx49590), .A0 (ram_131__6), .A1 (nx65580), .S0 (
             nx63632)) ;
    dffr reg_ram_130__6 (.Q (ram_130__6), .QB (\$dummy [1731]), .D (nx49600), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49601 (.Y (nx49600), .A0 (ram_130__6), .A1 (nx65580), .S0 (
             nx63636)) ;
    aoi22 ix61922 (.Y (nx61921), .A0 (ram_132__6), .A1 (nx64670), .B0 (
          ram_133__6), .B1 (nx64708)) ;
    dffr reg_ram_132__6 (.Q (ram_132__6), .QB (\$dummy [1732]), .D (nx49580), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49581 (.Y (nx49580), .A0 (ram_132__6), .A1 (nx65582), .S0 (
             nx63628)) ;
    dffr reg_ram_133__6 (.Q (ram_133__6), .QB (\$dummy [1733]), .D (nx49570), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49571 (.Y (nx49570), .A0 (ram_133__6), .A1 (nx65582), .S0 (
             nx63624)) ;
    aoi22 ix61930 (.Y (nx61929), .A0 (ram_135__6), .A1 (nx64746), .B0 (
          ram_134__6), .B1 (nx64784)) ;
    dffr reg_ram_135__6 (.Q (ram_135__6), .QB (\$dummy [1734]), .D (nx49550), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49551 (.Y (nx49550), .A0 (ram_135__6), .A1 (nx65582), .S0 (
             nx63616)) ;
    dffr reg_ram_134__6 (.Q (ram_134__6), .QB (\$dummy [1735]), .D (nx49560), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49561 (.Y (nx49560), .A0 (ram_134__6), .A1 (nx65582), .S0 (
             nx63620)) ;
    nand04 ix18473 (.Y (nx18472), .A0 (nx61938), .A1 (nx61946), .A2 (nx61954), .A3 (
           nx61962)) ;
    aoi22 ix61939 (.Y (nx61938), .A0 (ram_136__6), .A1 (nx64822), .B0 (
          ram_137__6), .B1 (nx64860)) ;
    dffr reg_ram_136__6 (.Q (ram_136__6), .QB (\$dummy [1736]), .D (nx49540), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49541 (.Y (nx49540), .A0 (ram_136__6), .A1 (nx65582), .S0 (
             nx63612)) ;
    dffr reg_ram_137__6 (.Q (ram_137__6), .QB (\$dummy [1737]), .D (nx49530), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49531 (.Y (nx49530), .A0 (ram_137__6), .A1 (nx65582), .S0 (
             nx63608)) ;
    aoi22 ix61947 (.Y (nx61946), .A0 (ram_139__6), .A1 (nx64898), .B0 (
          ram_138__6), .B1 (nx64936)) ;
    dffr reg_ram_139__6 (.Q (ram_139__6), .QB (\$dummy [1738]), .D (nx49510), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49511 (.Y (nx49510), .A0 (ram_139__6), .A1 (nx65582), .S0 (
             nx63600)) ;
    dffr reg_ram_138__6 (.Q (ram_138__6), .QB (\$dummy [1739]), .D (nx49520), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49521 (.Y (nx49520), .A0 (ram_138__6), .A1 (nx65584), .S0 (
             nx63604)) ;
    aoi22 ix61955 (.Y (nx61954), .A0 (ram_140__6), .A1 (nx64974), .B0 (
          ram_141__6), .B1 (nx65012)) ;
    dffr reg_ram_140__6 (.Q (ram_140__6), .QB (\$dummy [1740]), .D (nx49500), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49501 (.Y (nx49500), .A0 (ram_140__6), .A1 (nx65584), .S0 (
             nx63596)) ;
    dffr reg_ram_141__6 (.Q (ram_141__6), .QB (\$dummy [1741]), .D (nx49490), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49491 (.Y (nx49490), .A0 (ram_141__6), .A1 (nx65584), .S0 (
             nx63592)) ;
    aoi22 ix61963 (.Y (nx61962), .A0 (ram_143__6), .A1 (nx65050), .B0 (
          ram_142__6), .B1 (nx65088)) ;
    dffr reg_ram_143__6 (.Q (ram_143__6), .QB (\$dummy [1742]), .D (nx49470), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49471 (.Y (nx49470), .A0 (ram_143__6), .A1 (nx65584), .S0 (
             nx63584)) ;
    dffr reg_ram_142__6 (.Q (ram_142__6), .QB (\$dummy [1743]), .D (nx49480), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49481 (.Y (nx49480), .A0 (ram_142__6), .A1 (nx65584), .S0 (
             nx63588)) ;
    oai21 ix61971 (.Y (nx61970), .A0 (nx18388), .A1 (nx18310), .B0 (nx65218)) ;
    nand04 ix18389 (.Y (nx18388), .A0 (nx61973), .A1 (nx61981), .A2 (nx61989), .A3 (
           nx61997)) ;
    aoi22 ix61974 (.Y (nx61973), .A0 (ram_144__6), .A1 (nx64518), .B0 (
          ram_145__6), .B1 (nx64556)) ;
    dffr reg_ram_144__6 (.Q (ram_144__6), .QB (\$dummy [1744]), .D (nx49460), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49461 (.Y (nx49460), .A0 (ram_144__6), .A1 (nx65584), .S0 (
             nx63574)) ;
    dffr reg_ram_145__6 (.Q (ram_145__6), .QB (\$dummy [1745]), .D (nx49450), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49451 (.Y (nx49450), .A0 (ram_145__6), .A1 (nx65584), .S0 (
             nx63570)) ;
    aoi22 ix61982 (.Y (nx61981), .A0 (ram_147__6), .A1 (nx64594), .B0 (
          ram_146__6), .B1 (nx64632)) ;
    dffr reg_ram_147__6 (.Q (ram_147__6), .QB (\$dummy [1746]), .D (nx49430), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49431 (.Y (nx49430), .A0 (ram_147__6), .A1 (nx65586), .S0 (
             nx63562)) ;
    dffr reg_ram_146__6 (.Q (ram_146__6), .QB (\$dummy [1747]), .D (nx49440), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49441 (.Y (nx49440), .A0 (ram_146__6), .A1 (nx65586), .S0 (
             nx63566)) ;
    aoi22 ix61990 (.Y (nx61989), .A0 (ram_148__6), .A1 (nx64670), .B0 (
          ram_149__6), .B1 (nx64708)) ;
    dffr reg_ram_148__6 (.Q (ram_148__6), .QB (\$dummy [1748]), .D (nx49420), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49421 (.Y (nx49420), .A0 (ram_148__6), .A1 (nx65586), .S0 (
             nx63558)) ;
    dffr reg_ram_149__6 (.Q (ram_149__6), .QB (\$dummy [1749]), .D (nx49410), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49411 (.Y (nx49410), .A0 (ram_149__6), .A1 (nx65586), .S0 (
             nx63554)) ;
    aoi22 ix61998 (.Y (nx61997), .A0 (ram_151__6), .A1 (nx64746), .B0 (
          ram_150__6), .B1 (nx64784)) ;
    dffr reg_ram_151__6 (.Q (ram_151__6), .QB (\$dummy [1750]), .D (nx49390), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49391 (.Y (nx49390), .A0 (ram_151__6), .A1 (nx65586), .S0 (
             nx63546)) ;
    dffr reg_ram_150__6 (.Q (ram_150__6), .QB (\$dummy [1751]), .D (nx49400), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49401 (.Y (nx49400), .A0 (ram_150__6), .A1 (nx65586), .S0 (
             nx63550)) ;
    nand04 ix18311 (.Y (nx18310), .A0 (nx62006), .A1 (nx62014), .A2 (nx62022), .A3 (
           nx62030)) ;
    aoi22 ix62007 (.Y (nx62006), .A0 (ram_152__6), .A1 (nx64822), .B0 (
          ram_153__6), .B1 (nx64860)) ;
    dffr reg_ram_152__6 (.Q (ram_152__6), .QB (\$dummy [1752]), .D (nx49380), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49381 (.Y (nx49380), .A0 (ram_152__6), .A1 (nx65586), .S0 (
             nx63542)) ;
    dffr reg_ram_153__6 (.Q (ram_153__6), .QB (\$dummy [1753]), .D (nx49370), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49371 (.Y (nx49370), .A0 (ram_153__6), .A1 (nx65588), .S0 (
             nx63538)) ;
    aoi22 ix62015 (.Y (nx62014), .A0 (ram_155__6), .A1 (nx64898), .B0 (
          ram_154__6), .B1 (nx64936)) ;
    dffr reg_ram_155__6 (.Q (ram_155__6), .QB (\$dummy [1754]), .D (nx49350), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49351 (.Y (nx49350), .A0 (ram_155__6), .A1 (nx65588), .S0 (
             nx63530)) ;
    dffr reg_ram_154__6 (.Q (ram_154__6), .QB (\$dummy [1755]), .D (nx49360), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49361 (.Y (nx49360), .A0 (ram_154__6), .A1 (nx65588), .S0 (
             nx63534)) ;
    aoi22 ix62023 (.Y (nx62022), .A0 (ram_156__6), .A1 (nx64974), .B0 (
          ram_157__6), .B1 (nx65012)) ;
    dffr reg_ram_156__6 (.Q (ram_156__6), .QB (\$dummy [1756]), .D (nx49340), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49341 (.Y (nx49340), .A0 (ram_156__6), .A1 (nx65588), .S0 (
             nx63526)) ;
    dffr reg_ram_157__6 (.Q (ram_157__6), .QB (\$dummy [1757]), .D (nx49330), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49331 (.Y (nx49330), .A0 (ram_157__6), .A1 (nx65588), .S0 (
             nx63522)) ;
    aoi22 ix62031 (.Y (nx62030), .A0 (ram_159__6), .A1 (nx65050), .B0 (
          ram_158__6), .B1 (nx65088)) ;
    dffr reg_ram_159__6 (.Q (ram_159__6), .QB (\$dummy [1758]), .D (nx49310), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49311 (.Y (nx49310), .A0 (ram_159__6), .A1 (nx65588), .S0 (
             nx63514)) ;
    dffr reg_ram_158__6 (.Q (ram_158__6), .QB (\$dummy [1759]), .D (nx49320), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49321 (.Y (nx49320), .A0 (ram_158__6), .A1 (nx65588), .S0 (
             nx63518)) ;
    oai21 ix62039 (.Y (nx62038), .A0 (nx18224), .A1 (nx18146), .B0 (nx65222)) ;
    nand04 ix18225 (.Y (nx18224), .A0 (nx62041), .A1 (nx62049), .A2 (nx62057), .A3 (
           nx62065)) ;
    aoi22 ix62042 (.Y (nx62041), .A0 (ram_160__6), .A1 (nx64518), .B0 (
          ram_161__6), .B1 (nx64556)) ;
    dffr reg_ram_160__6 (.Q (ram_160__6), .QB (\$dummy [1760]), .D (nx49300), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49301 (.Y (nx49300), .A0 (ram_160__6), .A1 (nx65590), .S0 (
             nx63504)) ;
    dffr reg_ram_161__6 (.Q (ram_161__6), .QB (\$dummy [1761]), .D (nx49290), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49291 (.Y (nx49290), .A0 (ram_161__6), .A1 (nx65590), .S0 (
             nx63500)) ;
    aoi22 ix62050 (.Y (nx62049), .A0 (ram_163__6), .A1 (nx64594), .B0 (
          ram_162__6), .B1 (nx64632)) ;
    dffr reg_ram_163__6 (.Q (ram_163__6), .QB (\$dummy [1762]), .D (nx49270), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49271 (.Y (nx49270), .A0 (ram_163__6), .A1 (nx65590), .S0 (
             nx63492)) ;
    dffr reg_ram_162__6 (.Q (ram_162__6), .QB (\$dummy [1763]), .D (nx49280), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49281 (.Y (nx49280), .A0 (ram_162__6), .A1 (nx65590), .S0 (
             nx63496)) ;
    aoi22 ix62058 (.Y (nx62057), .A0 (ram_164__6), .A1 (nx64670), .B0 (
          ram_165__6), .B1 (nx64708)) ;
    dffr reg_ram_164__6 (.Q (ram_164__6), .QB (\$dummy [1764]), .D (nx49260), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49261 (.Y (nx49260), .A0 (ram_164__6), .A1 (nx65590), .S0 (
             nx63488)) ;
    dffr reg_ram_165__6 (.Q (ram_165__6), .QB (\$dummy [1765]), .D (nx49250), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49251 (.Y (nx49250), .A0 (ram_165__6), .A1 (nx65590), .S0 (
             nx63484)) ;
    aoi22 ix62066 (.Y (nx62065), .A0 (ram_167__6), .A1 (nx64746), .B0 (
          ram_166__6), .B1 (nx64784)) ;
    dffr reg_ram_167__6 (.Q (ram_167__6), .QB (\$dummy [1766]), .D (nx49230), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49231 (.Y (nx49230), .A0 (ram_167__6), .A1 (nx65590), .S0 (
             nx63476)) ;
    dffr reg_ram_166__6 (.Q (ram_166__6), .QB (\$dummy [1767]), .D (nx49240), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49241 (.Y (nx49240), .A0 (ram_166__6), .A1 (nx65592), .S0 (
             nx63480)) ;
    nand04 ix18147 (.Y (nx18146), .A0 (nx62074), .A1 (nx62082), .A2 (nx62090), .A3 (
           nx62098)) ;
    aoi22 ix62075 (.Y (nx62074), .A0 (ram_168__6), .A1 (nx64822), .B0 (
          ram_169__6), .B1 (nx64860)) ;
    dffr reg_ram_168__6 (.Q (ram_168__6), .QB (\$dummy [1768]), .D (nx49220), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49221 (.Y (nx49220), .A0 (ram_168__6), .A1 (nx65592), .S0 (
             nx63472)) ;
    dffr reg_ram_169__6 (.Q (ram_169__6), .QB (\$dummy [1769]), .D (nx49210), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49211 (.Y (nx49210), .A0 (ram_169__6), .A1 (nx65592), .S0 (
             nx63468)) ;
    aoi22 ix62083 (.Y (nx62082), .A0 (ram_171__6), .A1 (nx64898), .B0 (
          ram_170__6), .B1 (nx64936)) ;
    dffr reg_ram_171__6 (.Q (ram_171__6), .QB (\$dummy [1770]), .D (nx49190), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49191 (.Y (nx49190), .A0 (ram_171__6), .A1 (nx65592), .S0 (
             nx63460)) ;
    dffr reg_ram_170__6 (.Q (ram_170__6), .QB (\$dummy [1771]), .D (nx49200), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49201 (.Y (nx49200), .A0 (ram_170__6), .A1 (nx65592), .S0 (
             nx63464)) ;
    aoi22 ix62091 (.Y (nx62090), .A0 (ram_172__6), .A1 (nx64974), .B0 (
          ram_173__6), .B1 (nx65012)) ;
    dffr reg_ram_172__6 (.Q (ram_172__6), .QB (\$dummy [1772]), .D (nx49180), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49181 (.Y (nx49180), .A0 (ram_172__6), .A1 (nx65592), .S0 (
             nx63456)) ;
    dffr reg_ram_173__6 (.Q (ram_173__6), .QB (\$dummy [1773]), .D (nx49170), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49171 (.Y (nx49170), .A0 (ram_173__6), .A1 (nx65592), .S0 (
             nx63452)) ;
    aoi22 ix62099 (.Y (nx62098), .A0 (ram_175__6), .A1 (nx65050), .B0 (
          ram_174__6), .B1 (nx65088)) ;
    dffr reg_ram_175__6 (.Q (ram_175__6), .QB (\$dummy [1774]), .D (nx49150), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49151 (.Y (nx49150), .A0 (ram_175__6), .A1 (nx65594), .S0 (
             nx63444)) ;
    dffr reg_ram_174__6 (.Q (ram_174__6), .QB (\$dummy [1775]), .D (nx49160), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49161 (.Y (nx49160), .A0 (ram_174__6), .A1 (nx65594), .S0 (
             nx63448)) ;
    oai21 ix62107 (.Y (nx62106), .A0 (nx18062), .A1 (nx17984), .B0 (nx65226)) ;
    nand04 ix18063 (.Y (nx18062), .A0 (nx62109), .A1 (nx62117), .A2 (nx62125), .A3 (
           nx62133)) ;
    aoi22 ix62110 (.Y (nx62109), .A0 (ram_176__6), .A1 (nx64520), .B0 (
          ram_177__6), .B1 (nx64558)) ;
    dffr reg_ram_176__6 (.Q (ram_176__6), .QB (\$dummy [1776]), .D (nx49140), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49141 (.Y (nx49140), .A0 (ram_176__6), .A1 (nx65594), .S0 (
             nx63434)) ;
    dffr reg_ram_177__6 (.Q (ram_177__6), .QB (\$dummy [1777]), .D (nx49130), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49131 (.Y (nx49130), .A0 (ram_177__6), .A1 (nx65594), .S0 (
             nx63424)) ;
    aoi22 ix62118 (.Y (nx62117), .A0 (ram_179__6), .A1 (nx64596), .B0 (
          ram_178__6), .B1 (nx64634)) ;
    dffr reg_ram_179__6 (.Q (ram_179__6), .QB (\$dummy [1778]), .D (nx49110), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49111 (.Y (nx49110), .A0 (ram_179__6), .A1 (nx65594), .S0 (
             nx63404)) ;
    dffr reg_ram_178__6 (.Q (ram_178__6), .QB (\$dummy [1779]), .D (nx49120), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49121 (.Y (nx49120), .A0 (ram_178__6), .A1 (nx65594), .S0 (
             nx63414)) ;
    aoi22 ix62126 (.Y (nx62125), .A0 (ram_180__6), .A1 (nx64672), .B0 (
          ram_181__6), .B1 (nx64710)) ;
    dffr reg_ram_180__6 (.Q (ram_180__6), .QB (\$dummy [1780]), .D (nx49100), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49101 (.Y (nx49100), .A0 (ram_180__6), .A1 (nx65594), .S0 (
             nx63394)) ;
    dffr reg_ram_181__6 (.Q (ram_181__6), .QB (\$dummy [1781]), .D (nx49090), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49091 (.Y (nx49090), .A0 (ram_181__6), .A1 (nx65596), .S0 (
             nx63384)) ;
    aoi22 ix62134 (.Y (nx62133), .A0 (ram_183__6), .A1 (nx64748), .B0 (
          ram_182__6), .B1 (nx64786)) ;
    dffr reg_ram_183__6 (.Q (ram_183__6), .QB (\$dummy [1782]), .D (nx49070), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49071 (.Y (nx49070), .A0 (ram_183__6), .A1 (nx65596), .S0 (
             nx63364)) ;
    dffr reg_ram_182__6 (.Q (ram_182__6), .QB (\$dummy [1783]), .D (nx49080), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49081 (.Y (nx49080), .A0 (ram_182__6), .A1 (nx65596), .S0 (
             nx63374)) ;
    nand04 ix17985 (.Y (nx17984), .A0 (nx62142), .A1 (nx62150), .A2 (nx62158), .A3 (
           nx62166)) ;
    aoi22 ix62143 (.Y (nx62142), .A0 (ram_184__6), .A1 (nx64824), .B0 (
          ram_185__6), .B1 (nx64862)) ;
    dffr reg_ram_184__6 (.Q (ram_184__6), .QB (\$dummy [1784]), .D (nx49060), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49061 (.Y (nx49060), .A0 (ram_184__6), .A1 (nx65596), .S0 (
             nx63354)) ;
    dffr reg_ram_185__6 (.Q (ram_185__6), .QB (\$dummy [1785]), .D (nx49050), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49051 (.Y (nx49050), .A0 (ram_185__6), .A1 (nx65596), .S0 (
             nx63344)) ;
    aoi22 ix62151 (.Y (nx62150), .A0 (ram_187__6), .A1 (nx64900), .B0 (
          ram_186__6), .B1 (nx64938)) ;
    dffr reg_ram_187__6 (.Q (ram_187__6), .QB (\$dummy [1786]), .D (nx49030), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49031 (.Y (nx49030), .A0 (ram_187__6), .A1 (nx65596), .S0 (
             nx63324)) ;
    dffr reg_ram_186__6 (.Q (ram_186__6), .QB (\$dummy [1787]), .D (nx49040), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49041 (.Y (nx49040), .A0 (ram_186__6), .A1 (nx65596), .S0 (
             nx63334)) ;
    aoi22 ix62159 (.Y (nx62158), .A0 (ram_188__6), .A1 (nx64976), .B0 (
          ram_189__6), .B1 (nx65014)) ;
    dffr reg_ram_188__6 (.Q (ram_188__6), .QB (\$dummy [1788]), .D (nx49020), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49021 (.Y (nx49020), .A0 (ram_188__6), .A1 (nx65598), .S0 (
             nx63314)) ;
    dffr reg_ram_189__6 (.Q (ram_189__6), .QB (\$dummy [1789]), .D (nx49010), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49011 (.Y (nx49010), .A0 (ram_189__6), .A1 (nx65598), .S0 (
             nx63304)) ;
    aoi22 ix62167 (.Y (nx62166), .A0 (ram_191__6), .A1 (nx65052), .B0 (
          ram_190__6), .B1 (nx65090)) ;
    dffr reg_ram_191__6 (.Q (ram_191__6), .QB (\$dummy [1790]), .D (nx48990), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix48991 (.Y (nx48990), .A0 (ram_191__6), .A1 (nx65598), .S0 (
             nx63284)) ;
    dffr reg_ram_190__6 (.Q (ram_190__6), .QB (\$dummy [1791]), .D (nx49000), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix49001 (.Y (nx49000), .A0 (ram_190__6), .A1 (nx65598), .S0 (
             nx63294)) ;
    or04 ix23151 (.Y (dataout[7]), .A0 (nx23146), .A1 (nx22492), .A2 (nx21836), 
         .A3 (nx21182)) ;
    nand04 ix23147 (.Y (nx23146), .A0 (nx62176), .A1 (nx62244), .A2 (nx62312), .A3 (
           nx62380)) ;
    oai21 ix62177 (.Y (nx62176), .A0 (nx23136), .A1 (nx23058), .B0 (nx66120)) ;
    nand04 ix23137 (.Y (nx23136), .A0 (nx62179), .A1 (nx62187), .A2 (nx62195), .A3 (
           nx62203)) ;
    aoi22 ix62180 (.Y (nx62179), .A0 (ram_240__7), .A1 (nx64520), .B0 (
          ram_241__7), .B1 (nx64558)) ;
    dffr reg_ram_240__7 (.Q (ram_240__7), .QB (\$dummy [1792]), .D (nx54100), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix54101 (.Y (nx54100), .A0 (ram_240__7), .A1 (nx65450), .S0 (
             nx64416)) ;
    dffr reg_ram_241__7 (.Q (ram_241__7), .QB (\$dummy [1793]), .D (nx54090), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix54091 (.Y (nx54090), .A0 (ram_241__7), .A1 (nx65450), .S0 (
             nx64412)) ;
    aoi22 ix62188 (.Y (nx62187), .A0 (ram_243__7), .A1 (nx64596), .B0 (
          ram_242__7), .B1 (nx64634)) ;
    dffr reg_ram_243__7 (.Q (ram_243__7), .QB (\$dummy [1794]), .D (nx54070), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix54071 (.Y (nx54070), .A0 (ram_243__7), .A1 (nx65450), .S0 (
             nx64404)) ;
    dffr reg_ram_242__7 (.Q (ram_242__7), .QB (\$dummy [1795]), .D (nx54080), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix54081 (.Y (nx54080), .A0 (ram_242__7), .A1 (nx65450), .S0 (
             nx64408)) ;
    aoi22 ix62196 (.Y (nx62195), .A0 (ram_244__7), .A1 (nx64672), .B0 (
          ram_245__7), .B1 (nx64710)) ;
    dffr reg_ram_244__7 (.Q (ram_244__7), .QB (\$dummy [1796]), .D (nx54060), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix54061 (.Y (nx54060), .A0 (ram_244__7), .A1 (nx65450), .S0 (
             nx64400)) ;
    dffr reg_ram_245__7 (.Q (ram_245__7), .QB (\$dummy [1797]), .D (nx54050), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix54051 (.Y (nx54050), .A0 (ram_245__7), .A1 (nx65450), .S0 (
             nx64396)) ;
    aoi22 ix62204 (.Y (nx62203), .A0 (ram_247__7), .A1 (nx64748), .B0 (
          ram_246__7), .B1 (nx64786)) ;
    dffr reg_ram_247__7 (.Q (ram_247__7), .QB (\$dummy [1798]), .D (nx54030), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix54031 (.Y (nx54030), .A0 (ram_247__7), .A1 (nx65450), .S0 (
             nx64388)) ;
    dffr reg_ram_246__7 (.Q (ram_246__7), .QB (\$dummy [1799]), .D (nx54040), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix54041 (.Y (nx54040), .A0 (ram_246__7), .A1 (nx65452), .S0 (
             nx64392)) ;
    nand04 ix23059 (.Y (nx23058), .A0 (nx62212), .A1 (nx62220), .A2 (nx62228), .A3 (
           nx62236)) ;
    aoi22 ix62213 (.Y (nx62212), .A0 (ram_248__7), .A1 (nx64824), .B0 (
          ram_249__7), .B1 (nx64862)) ;
    dffr reg_ram_248__7 (.Q (ram_248__7), .QB (\$dummy [1800]), .D (nx54020), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix54021 (.Y (nx54020), .A0 (ram_248__7), .A1 (nx65452), .S0 (
             nx64384)) ;
    dffr reg_ram_249__7 (.Q (ram_249__7), .QB (\$dummy [1801]), .D (nx54010), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix54011 (.Y (nx54010), .A0 (ram_249__7), .A1 (nx65452), .S0 (
             nx64380)) ;
    aoi22 ix62221 (.Y (nx62220), .A0 (ram_251__7), .A1 (nx64900), .B0 (
          ram_250__7), .B1 (nx64938)) ;
    dffr reg_ram_251__7 (.Q (ram_251__7), .QB (\$dummy [1802]), .D (nx53990), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53991 (.Y (nx53990), .A0 (ram_251__7), .A1 (nx65452), .S0 (
             nx64372)) ;
    dffr reg_ram_250__7 (.Q (ram_250__7), .QB (\$dummy [1803]), .D (nx54000), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix54001 (.Y (nx54000), .A0 (ram_250__7), .A1 (nx65452), .S0 (
             nx64376)) ;
    aoi22 ix62229 (.Y (nx62228), .A0 (ram_252__7), .A1 (nx64976), .B0 (
          ram_253__7), .B1 (nx65014)) ;
    dffr reg_ram_252__7 (.Q (ram_252__7), .QB (\$dummy [1804]), .D (nx53980), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53981 (.Y (nx53980), .A0 (ram_252__7), .A1 (nx65452), .S0 (
             nx64368)) ;
    dffr reg_ram_253__7 (.Q (ram_253__7), .QB (\$dummy [1805]), .D (nx53970), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53971 (.Y (nx53970), .A0 (ram_253__7), .A1 (nx65452), .S0 (
             nx64364)) ;
    aoi22 ix62237 (.Y (nx62236), .A0 (ram_255__7), .A1 (nx65052), .B0 (
          ram_254__7), .B1 (nx65090)) ;
    dffr reg_ram_255__7 (.Q (ram_255__7), .QB (\$dummy [1806]), .D (nx53950), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53951 (.Y (nx53950), .A0 (ram_255__7), .A1 (nx65454), .S0 (
             nx64356)) ;
    dffr reg_ram_254__7 (.Q (ram_254__7), .QB (\$dummy [1807]), .D (nx53960), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53961 (.Y (nx53960), .A0 (ram_254__7), .A1 (nx65454), .S0 (
             nx64360)) ;
    oai21 ix62245 (.Y (nx62244), .A0 (nx22974), .A1 (nx22896), .B0 (nx66124)) ;
    nand04 ix22975 (.Y (nx22974), .A0 (nx62247), .A1 (nx62255), .A2 (nx62263), .A3 (
           nx62271)) ;
    aoi22 ix62248 (.Y (nx62247), .A0 (ram_224__7), .A1 (nx64520), .B0 (
          ram_225__7), .B1 (nx64558)) ;
    dffr reg_ram_224__7 (.Q (ram_224__7), .QB (\$dummy [1808]), .D (nx53940), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53941 (.Y (nx53940), .A0 (ram_224__7), .A1 (nx65454), .S0 (
             nx64346)) ;
    dffr reg_ram_225__7 (.Q (ram_225__7), .QB (\$dummy [1809]), .D (nx53930), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53931 (.Y (nx53930), .A0 (ram_225__7), .A1 (nx65454), .S0 (
             nx64342)) ;
    aoi22 ix62256 (.Y (nx62255), .A0 (ram_227__7), .A1 (nx64596), .B0 (
          ram_226__7), .B1 (nx64634)) ;
    dffr reg_ram_227__7 (.Q (ram_227__7), .QB (\$dummy [1810]), .D (nx53910), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53911 (.Y (nx53910), .A0 (ram_227__7), .A1 (nx65454), .S0 (
             nx64334)) ;
    dffr reg_ram_226__7 (.Q (ram_226__7), .QB (\$dummy [1811]), .D (nx53920), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53921 (.Y (nx53920), .A0 (ram_226__7), .A1 (nx65454), .S0 (
             nx64338)) ;
    aoi22 ix62264 (.Y (nx62263), .A0 (ram_228__7), .A1 (nx64672), .B0 (
          ram_229__7), .B1 (nx64710)) ;
    dffr reg_ram_228__7 (.Q (ram_228__7), .QB (\$dummy [1812]), .D (nx53900), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53901 (.Y (nx53900), .A0 (ram_228__7), .A1 (nx65454), .S0 (
             nx64330)) ;
    dffr reg_ram_229__7 (.Q (ram_229__7), .QB (\$dummy [1813]), .D (nx53890), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53891 (.Y (nx53890), .A0 (ram_229__7), .A1 (nx65456), .S0 (
             nx64326)) ;
    aoi22 ix62272 (.Y (nx62271), .A0 (ram_231__7), .A1 (nx64748), .B0 (
          ram_230__7), .B1 (nx64786)) ;
    dffr reg_ram_231__7 (.Q (ram_231__7), .QB (\$dummy [1814]), .D (nx53870), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53871 (.Y (nx53870), .A0 (ram_231__7), .A1 (nx65456), .S0 (
             nx64318)) ;
    dffr reg_ram_230__7 (.Q (ram_230__7), .QB (\$dummy [1815]), .D (nx53880), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53881 (.Y (nx53880), .A0 (ram_230__7), .A1 (nx65456), .S0 (
             nx64322)) ;
    nand04 ix22897 (.Y (nx22896), .A0 (nx62280), .A1 (nx62288), .A2 (nx62296), .A3 (
           nx62304)) ;
    aoi22 ix62281 (.Y (nx62280), .A0 (ram_232__7), .A1 (nx64824), .B0 (
          ram_233__7), .B1 (nx64862)) ;
    dffr reg_ram_232__7 (.Q (ram_232__7), .QB (\$dummy [1816]), .D (nx53860), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53861 (.Y (nx53860), .A0 (ram_232__7), .A1 (nx65456), .S0 (
             nx64314)) ;
    dffr reg_ram_233__7 (.Q (ram_233__7), .QB (\$dummy [1817]), .D (nx53850), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53851 (.Y (nx53850), .A0 (ram_233__7), .A1 (nx65456), .S0 (
             nx64310)) ;
    aoi22 ix62289 (.Y (nx62288), .A0 (ram_235__7), .A1 (nx64900), .B0 (
          ram_234__7), .B1 (nx64938)) ;
    dffr reg_ram_235__7 (.Q (ram_235__7), .QB (\$dummy [1818]), .D (nx53830), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53831 (.Y (nx53830), .A0 (ram_235__7), .A1 (nx65456), .S0 (
             nx64302)) ;
    dffr reg_ram_234__7 (.Q (ram_234__7), .QB (\$dummy [1819]), .D (nx53840), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53841 (.Y (nx53840), .A0 (ram_234__7), .A1 (nx65456), .S0 (
             nx64306)) ;
    aoi22 ix62297 (.Y (nx62296), .A0 (ram_236__7), .A1 (nx64976), .B0 (
          ram_237__7), .B1 (nx65014)) ;
    dffr reg_ram_236__7 (.Q (ram_236__7), .QB (\$dummy [1820]), .D (nx53820), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53821 (.Y (nx53820), .A0 (ram_236__7), .A1 (nx65458), .S0 (
             nx64298)) ;
    dffr reg_ram_237__7 (.Q (ram_237__7), .QB (\$dummy [1821]), .D (nx53810), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53811 (.Y (nx53810), .A0 (ram_237__7), .A1 (nx65458), .S0 (
             nx64294)) ;
    aoi22 ix62305 (.Y (nx62304), .A0 (ram_239__7), .A1 (nx65052), .B0 (
          ram_238__7), .B1 (nx65090)) ;
    dffr reg_ram_239__7 (.Q (ram_239__7), .QB (\$dummy [1822]), .D (nx53790), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53791 (.Y (nx53790), .A0 (ram_239__7), .A1 (nx65458), .S0 (
             nx64286)) ;
    dffr reg_ram_238__7 (.Q (ram_238__7), .QB (\$dummy [1823]), .D (nx53800), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53801 (.Y (nx53800), .A0 (ram_238__7), .A1 (nx65458), .S0 (
             nx64290)) ;
    oai21 ix62313 (.Y (nx62312), .A0 (nx22810), .A1 (nx22732), .B0 (nx66128)) ;
    nand04 ix22811 (.Y (nx22810), .A0 (nx62315), .A1 (nx62323), .A2 (nx62331), .A3 (
           nx62339)) ;
    aoi22 ix62316 (.Y (nx62315), .A0 (ram_208__7), .A1 (nx64520), .B0 (
          ram_209__7), .B1 (nx64558)) ;
    dffr reg_ram_208__7 (.Q (ram_208__7), .QB (\$dummy [1824]), .D (nx53780), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53781 (.Y (nx53780), .A0 (ram_208__7), .A1 (nx65458), .S0 (
             nx64276)) ;
    dffr reg_ram_209__7 (.Q (ram_209__7), .QB (\$dummy [1825]), .D (nx53770), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53771 (.Y (nx53770), .A0 (ram_209__7), .A1 (nx65458), .S0 (
             nx64272)) ;
    aoi22 ix62324 (.Y (nx62323), .A0 (ram_211__7), .A1 (nx64596), .B0 (
          ram_210__7), .B1 (nx64634)) ;
    dffr reg_ram_211__7 (.Q (ram_211__7), .QB (\$dummy [1826]), .D (nx53750), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53751 (.Y (nx53750), .A0 (ram_211__7), .A1 (nx65458), .S0 (
             nx64264)) ;
    dffr reg_ram_210__7 (.Q (ram_210__7), .QB (\$dummy [1827]), .D (nx53760), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53761 (.Y (nx53760), .A0 (ram_210__7), .A1 (nx65460), .S0 (
             nx64268)) ;
    aoi22 ix62332 (.Y (nx62331), .A0 (ram_212__7), .A1 (nx64672), .B0 (
          ram_213__7), .B1 (nx64710)) ;
    dffr reg_ram_212__7 (.Q (ram_212__7), .QB (\$dummy [1828]), .D (nx53740), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53741 (.Y (nx53740), .A0 (ram_212__7), .A1 (nx65460), .S0 (
             nx64260)) ;
    dffr reg_ram_213__7 (.Q (ram_213__7), .QB (\$dummy [1829]), .D (nx53730), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53731 (.Y (nx53730), .A0 (ram_213__7), .A1 (nx65460), .S0 (
             nx64256)) ;
    aoi22 ix62340 (.Y (nx62339), .A0 (ram_215__7), .A1 (nx64748), .B0 (
          ram_214__7), .B1 (nx64786)) ;
    dffr reg_ram_215__7 (.Q (ram_215__7), .QB (\$dummy [1830]), .D (nx53710), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53711 (.Y (nx53710), .A0 (ram_215__7), .A1 (nx65460), .S0 (
             nx64248)) ;
    dffr reg_ram_214__7 (.Q (ram_214__7), .QB (\$dummy [1831]), .D (nx53720), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53721 (.Y (nx53720), .A0 (ram_214__7), .A1 (nx65460), .S0 (
             nx64252)) ;
    nand04 ix22733 (.Y (nx22732), .A0 (nx62348), .A1 (nx62356), .A2 (nx62364), .A3 (
           nx62372)) ;
    aoi22 ix62349 (.Y (nx62348), .A0 (ram_216__7), .A1 (nx64824), .B0 (
          ram_217__7), .B1 (nx64862)) ;
    dffr reg_ram_216__7 (.Q (ram_216__7), .QB (\$dummy [1832]), .D (nx53700), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53701 (.Y (nx53700), .A0 (ram_216__7), .A1 (nx65460), .S0 (
             nx64244)) ;
    dffr reg_ram_217__7 (.Q (ram_217__7), .QB (\$dummy [1833]), .D (nx53690), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53691 (.Y (nx53690), .A0 (ram_217__7), .A1 (nx65460), .S0 (
             nx64240)) ;
    aoi22 ix62357 (.Y (nx62356), .A0 (ram_219__7), .A1 (nx64900), .B0 (
          ram_218__7), .B1 (nx64938)) ;
    dffr reg_ram_219__7 (.Q (ram_219__7), .QB (\$dummy [1834]), .D (nx53670), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53671 (.Y (nx53670), .A0 (ram_219__7), .A1 (nx65462), .S0 (
             nx64232)) ;
    dffr reg_ram_218__7 (.Q (ram_218__7), .QB (\$dummy [1835]), .D (nx53680), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53681 (.Y (nx53680), .A0 (ram_218__7), .A1 (nx65462), .S0 (
             nx64236)) ;
    aoi22 ix62365 (.Y (nx62364), .A0 (ram_220__7), .A1 (nx64976), .B0 (
          ram_221__7), .B1 (nx65014)) ;
    dffr reg_ram_220__7 (.Q (ram_220__7), .QB (\$dummy [1836]), .D (nx53660), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53661 (.Y (nx53660), .A0 (ram_220__7), .A1 (nx65462), .S0 (
             nx64228)) ;
    dffr reg_ram_221__7 (.Q (ram_221__7), .QB (\$dummy [1837]), .D (nx53650), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53651 (.Y (nx53650), .A0 (ram_221__7), .A1 (nx65462), .S0 (
             nx64224)) ;
    aoi22 ix62373 (.Y (nx62372), .A0 (ram_223__7), .A1 (nx65052), .B0 (
          ram_222__7), .B1 (nx65090)) ;
    dffr reg_ram_223__7 (.Q (ram_223__7), .QB (\$dummy [1838]), .D (nx53630), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53631 (.Y (nx53630), .A0 (ram_223__7), .A1 (nx65462), .S0 (
             nx64216)) ;
    dffr reg_ram_222__7 (.Q (ram_222__7), .QB (\$dummy [1839]), .D (nx53640), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53641 (.Y (nx53640), .A0 (ram_222__7), .A1 (nx65462), .S0 (
             nx64220)) ;
    oai21 ix62381 (.Y (nx62380), .A0 (nx22648), .A1 (nx22570), .B0 (nx66132)) ;
    nand04 ix22649 (.Y (nx22648), .A0 (nx62383), .A1 (nx62391), .A2 (nx62399), .A3 (
           nx62407)) ;
    aoi22 ix62384 (.Y (nx62383), .A0 (ram_192__7), .A1 (nx64520), .B0 (
          ram_193__7), .B1 (nx64558)) ;
    dffr reg_ram_192__7 (.Q (ram_192__7), .QB (\$dummy [1840]), .D (nx53620), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53621 (.Y (nx53620), .A0 (ram_192__7), .A1 (nx65462), .S0 (
             nx64206)) ;
    dffr reg_ram_193__7 (.Q (ram_193__7), .QB (\$dummy [1841]), .D (nx53610), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53611 (.Y (nx53610), .A0 (ram_193__7), .A1 (nx65464), .S0 (
             nx64202)) ;
    aoi22 ix62392 (.Y (nx62391), .A0 (ram_195__7), .A1 (nx64596), .B0 (
          ram_194__7), .B1 (nx64634)) ;
    dffr reg_ram_195__7 (.Q (ram_195__7), .QB (\$dummy [1842]), .D (nx53590), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53591 (.Y (nx53590), .A0 (ram_195__7), .A1 (nx65464), .S0 (
             nx64194)) ;
    dffr reg_ram_194__7 (.Q (ram_194__7), .QB (\$dummy [1843]), .D (nx53600), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53601 (.Y (nx53600), .A0 (ram_194__7), .A1 (nx65464), .S0 (
             nx64198)) ;
    aoi22 ix62400 (.Y (nx62399), .A0 (ram_196__7), .A1 (nx64672), .B0 (
          ram_197__7), .B1 (nx64710)) ;
    dffr reg_ram_196__7 (.Q (ram_196__7), .QB (\$dummy [1844]), .D (nx53580), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53581 (.Y (nx53580), .A0 (ram_196__7), .A1 (nx65464), .S0 (
             nx64190)) ;
    dffr reg_ram_197__7 (.Q (ram_197__7), .QB (\$dummy [1845]), .D (nx53570), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53571 (.Y (nx53570), .A0 (ram_197__7), .A1 (nx65464), .S0 (
             nx64186)) ;
    aoi22 ix62408 (.Y (nx62407), .A0 (ram_199__7), .A1 (nx64748), .B0 (
          ram_198__7), .B1 (nx64786)) ;
    dffr reg_ram_199__7 (.Q (ram_199__7), .QB (\$dummy [1846]), .D (nx53550), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53551 (.Y (nx53550), .A0 (ram_199__7), .A1 (nx65464), .S0 (
             nx64178)) ;
    dffr reg_ram_198__7 (.Q (ram_198__7), .QB (\$dummy [1847]), .D (nx53560), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53561 (.Y (nx53560), .A0 (ram_198__7), .A1 (nx65464), .S0 (
             nx64182)) ;
    nand04 ix22571 (.Y (nx22570), .A0 (nx62416), .A1 (nx62424), .A2 (nx62432), .A3 (
           nx62440)) ;
    aoi22 ix62417 (.Y (nx62416), .A0 (ram_200__7), .A1 (nx64824), .B0 (
          ram_201__7), .B1 (nx64862)) ;
    dffr reg_ram_200__7 (.Q (ram_200__7), .QB (\$dummy [1848]), .D (nx53540), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53541 (.Y (nx53540), .A0 (ram_200__7), .A1 (nx65466), .S0 (
             nx64174)) ;
    dffr reg_ram_201__7 (.Q (ram_201__7), .QB (\$dummy [1849]), .D (nx53530), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53531 (.Y (nx53530), .A0 (ram_201__7), .A1 (nx65466), .S0 (
             nx64170)) ;
    aoi22 ix62425 (.Y (nx62424), .A0 (ram_203__7), .A1 (nx64900), .B0 (
          ram_202__7), .B1 (nx64938)) ;
    dffr reg_ram_203__7 (.Q (ram_203__7), .QB (\$dummy [1850]), .D (nx53510), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53511 (.Y (nx53510), .A0 (ram_203__7), .A1 (nx65466), .S0 (
             nx64162)) ;
    dffr reg_ram_202__7 (.Q (ram_202__7), .QB (\$dummy [1851]), .D (nx53520), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53521 (.Y (nx53520), .A0 (ram_202__7), .A1 (nx65466), .S0 (
             nx64166)) ;
    aoi22 ix62433 (.Y (nx62432), .A0 (ram_204__7), .A1 (nx64976), .B0 (
          ram_205__7), .B1 (nx65014)) ;
    dffr reg_ram_204__7 (.Q (ram_204__7), .QB (\$dummy [1852]), .D (nx53500), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53501 (.Y (nx53500), .A0 (ram_204__7), .A1 (nx65466), .S0 (
             nx64158)) ;
    dffr reg_ram_205__7 (.Q (ram_205__7), .QB (\$dummy [1853]), .D (nx53490), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53491 (.Y (nx53490), .A0 (ram_205__7), .A1 (nx65466), .S0 (
             nx64154)) ;
    aoi22 ix62441 (.Y (nx62440), .A0 (ram_207__7), .A1 (nx65052), .B0 (
          ram_206__7), .B1 (nx65090)) ;
    dffr reg_ram_207__7 (.Q (ram_207__7), .QB (\$dummy [1854]), .D (nx53470), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53471 (.Y (nx53470), .A0 (ram_207__7), .A1 (nx65466), .S0 (
             nx64146)) ;
    dffr reg_ram_206__7 (.Q (ram_206__7), .QB (\$dummy [1855]), .D (nx53480), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53481 (.Y (nx53480), .A0 (ram_206__7), .A1 (nx65468), .S0 (
             nx64150)) ;
    nand04 ix22493 (.Y (nx22492), .A0 (nx62449), .A1 (nx62517), .A2 (nx62585), .A3 (
           nx62653)) ;
    oai21 ix62450 (.Y (nx62449), .A0 (nx22482), .A1 (nx22404), .B0 (nx66136)) ;
    nand04 ix22483 (.Y (nx22482), .A0 (nx62452), .A1 (nx62460), .A2 (nx62468), .A3 (
           nx62476)) ;
    aoi22 ix62453 (.Y (nx62452), .A0 (ram_80__7), .A1 (nx64520), .B0 (ram_81__7)
          , .B1 (nx64558)) ;
    dffr reg_ram_80__7 (.Q (ram_80__7), .QB (\$dummy [1856]), .D (nx53460), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53461 (.Y (nx53460), .A0 (ram_80__7), .A1 (nx65468), .S0 (nx64136
             )) ;
    dffr reg_ram_81__7 (.Q (ram_81__7), .QB (\$dummy [1857]), .D (nx53450), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53451 (.Y (nx53450), .A0 (ram_81__7), .A1 (nx65468), .S0 (nx64132
             )) ;
    aoi22 ix62461 (.Y (nx62460), .A0 (ram_83__7), .A1 (nx64596), .B0 (ram_82__7)
          , .B1 (nx64634)) ;
    dffr reg_ram_83__7 (.Q (ram_83__7), .QB (\$dummy [1858]), .D (nx53430), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53431 (.Y (nx53430), .A0 (ram_83__7), .A1 (nx65468), .S0 (nx64124
             )) ;
    dffr reg_ram_82__7 (.Q (ram_82__7), .QB (\$dummy [1859]), .D (nx53440), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53441 (.Y (nx53440), .A0 (ram_82__7), .A1 (nx65468), .S0 (nx64128
             )) ;
    aoi22 ix62469 (.Y (nx62468), .A0 (ram_84__7), .A1 (nx64672), .B0 (ram_85__7)
          , .B1 (nx64710)) ;
    dffr reg_ram_84__7 (.Q (ram_84__7), .QB (\$dummy [1860]), .D (nx53420), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53421 (.Y (nx53420), .A0 (ram_84__7), .A1 (nx65468), .S0 (nx64120
             )) ;
    dffr reg_ram_85__7 (.Q (ram_85__7), .QB (\$dummy [1861]), .D (nx53410), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53411 (.Y (nx53410), .A0 (ram_85__7), .A1 (nx65468), .S0 (nx64116
             )) ;
    aoi22 ix62477 (.Y (nx62476), .A0 (ram_87__7), .A1 (nx64748), .B0 (ram_86__7)
          , .B1 (nx64786)) ;
    dffr reg_ram_87__7 (.Q (ram_87__7), .QB (\$dummy [1862]), .D (nx53390), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53391 (.Y (nx53390), .A0 (ram_87__7), .A1 (nx65470), .S0 (nx64108
             )) ;
    dffr reg_ram_86__7 (.Q (ram_86__7), .QB (\$dummy [1863]), .D (nx53400), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53401 (.Y (nx53400), .A0 (ram_86__7), .A1 (nx65470), .S0 (nx64112
             )) ;
    nand04 ix22405 (.Y (nx22404), .A0 (nx62485), .A1 (nx62493), .A2 (nx62501), .A3 (
           nx62509)) ;
    aoi22 ix62486 (.Y (nx62485), .A0 (ram_88__7), .A1 (nx64824), .B0 (ram_89__7)
          , .B1 (nx64862)) ;
    dffr reg_ram_88__7 (.Q (ram_88__7), .QB (\$dummy [1864]), .D (nx53380), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53381 (.Y (nx53380), .A0 (ram_88__7), .A1 (nx65470), .S0 (nx64104
             )) ;
    dffr reg_ram_89__7 (.Q (ram_89__7), .QB (\$dummy [1865]), .D (nx53370), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53371 (.Y (nx53370), .A0 (ram_89__7), .A1 (nx65470), .S0 (nx64100
             )) ;
    aoi22 ix62494 (.Y (nx62493), .A0 (ram_91__7), .A1 (nx64900), .B0 (ram_90__7)
          , .B1 (nx64938)) ;
    dffr reg_ram_91__7 (.Q (ram_91__7), .QB (\$dummy [1866]), .D (nx53350), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53351 (.Y (nx53350), .A0 (ram_91__7), .A1 (nx65470), .S0 (nx64092
             )) ;
    dffr reg_ram_90__7 (.Q (ram_90__7), .QB (\$dummy [1867]), .D (nx53360), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53361 (.Y (nx53360), .A0 (ram_90__7), .A1 (nx65470), .S0 (nx64096
             )) ;
    aoi22 ix62502 (.Y (nx62501), .A0 (ram_92__7), .A1 (nx64976), .B0 (ram_93__7)
          , .B1 (nx65014)) ;
    dffr reg_ram_92__7 (.Q (ram_92__7), .QB (\$dummy [1868]), .D (nx53340), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53341 (.Y (nx53340), .A0 (ram_92__7), .A1 (nx65470), .S0 (nx64088
             )) ;
    dffr reg_ram_93__7 (.Q (ram_93__7), .QB (\$dummy [1869]), .D (nx53330), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53331 (.Y (nx53330), .A0 (ram_93__7), .A1 (nx65472), .S0 (nx64084
             )) ;
    aoi22 ix62510 (.Y (nx62509), .A0 (ram_95__7), .A1 (nx65052), .B0 (ram_94__7)
          , .B1 (nx65090)) ;
    dffr reg_ram_95__7 (.Q (ram_95__7), .QB (\$dummy [1870]), .D (nx53310), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53311 (.Y (nx53310), .A0 (ram_95__7), .A1 (nx65472), .S0 (nx64076
             )) ;
    dffr reg_ram_94__7 (.Q (ram_94__7), .QB (\$dummy [1871]), .D (nx53320), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53321 (.Y (nx53320), .A0 (ram_94__7), .A1 (nx65472), .S0 (nx64080
             )) ;
    oai21 ix62518 (.Y (nx62517), .A0 (nx22320), .A1 (nx22242), .B0 (nx66140)) ;
    nand04 ix22321 (.Y (nx22320), .A0 (nx62520), .A1 (nx62528), .A2 (nx62536), .A3 (
           nx62544)) ;
    aoi22 ix62521 (.Y (nx62520), .A0 (ram_64__7), .A1 (nx64520), .B0 (ram_65__7)
          , .B1 (nx64558)) ;
    dffr reg_ram_64__7 (.Q (ram_64__7), .QB (\$dummy [1872]), .D (nx53300), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53301 (.Y (nx53300), .A0 (ram_64__7), .A1 (nx65472), .S0 (nx64066
             )) ;
    dffr reg_ram_65__7 (.Q (ram_65__7), .QB (\$dummy [1873]), .D (nx53290), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53291 (.Y (nx53290), .A0 (ram_65__7), .A1 (nx65472), .S0 (nx64062
             )) ;
    aoi22 ix62529 (.Y (nx62528), .A0 (ram_67__7), .A1 (nx64596), .B0 (ram_66__7)
          , .B1 (nx64634)) ;
    dffr reg_ram_67__7 (.Q (ram_67__7), .QB (\$dummy [1874]), .D (nx53270), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53271 (.Y (nx53270), .A0 (ram_67__7), .A1 (nx65472), .S0 (nx64054
             )) ;
    dffr reg_ram_66__7 (.Q (ram_66__7), .QB (\$dummy [1875]), .D (nx53280), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53281 (.Y (nx53280), .A0 (ram_66__7), .A1 (nx65472), .S0 (nx64058
             )) ;
    aoi22 ix62537 (.Y (nx62536), .A0 (ram_68__7), .A1 (nx64672), .B0 (ram_69__7)
          , .B1 (nx64710)) ;
    dffr reg_ram_68__7 (.Q (ram_68__7), .QB (\$dummy [1876]), .D (nx53260), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53261 (.Y (nx53260), .A0 (ram_68__7), .A1 (nx65474), .S0 (nx64050
             )) ;
    dffr reg_ram_69__7 (.Q (ram_69__7), .QB (\$dummy [1877]), .D (nx53250), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53251 (.Y (nx53250), .A0 (ram_69__7), .A1 (nx65474), .S0 (nx64046
             )) ;
    aoi22 ix62545 (.Y (nx62544), .A0 (ram_71__7), .A1 (nx64748), .B0 (ram_70__7)
          , .B1 (nx64786)) ;
    dffr reg_ram_71__7 (.Q (ram_71__7), .QB (\$dummy [1878]), .D (nx53230), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53231 (.Y (nx53230), .A0 (ram_71__7), .A1 (nx65474), .S0 (nx64038
             )) ;
    dffr reg_ram_70__7 (.Q (ram_70__7), .QB (\$dummy [1879]), .D (nx53240), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53241 (.Y (nx53240), .A0 (ram_70__7), .A1 (nx65474), .S0 (nx64042
             )) ;
    nand04 ix22243 (.Y (nx22242), .A0 (nx62553), .A1 (nx62561), .A2 (nx62569), .A3 (
           nx62577)) ;
    aoi22 ix62554 (.Y (nx62553), .A0 (ram_72__7), .A1 (nx64824), .B0 (ram_73__7)
          , .B1 (nx64862)) ;
    dffr reg_ram_72__7 (.Q (ram_72__7), .QB (\$dummy [1880]), .D (nx53220), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53221 (.Y (nx53220), .A0 (ram_72__7), .A1 (nx65474), .S0 (nx64034
             )) ;
    dffr reg_ram_73__7 (.Q (ram_73__7), .QB (\$dummy [1881]), .D (nx53210), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53211 (.Y (nx53210), .A0 (ram_73__7), .A1 (nx65474), .S0 (nx64030
             )) ;
    aoi22 ix62562 (.Y (nx62561), .A0 (ram_75__7), .A1 (nx64900), .B0 (ram_74__7)
          , .B1 (nx64938)) ;
    dffr reg_ram_75__7 (.Q (ram_75__7), .QB (\$dummy [1882]), .D (nx53190), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53191 (.Y (nx53190), .A0 (ram_75__7), .A1 (nx65474), .S0 (nx64022
             )) ;
    dffr reg_ram_74__7 (.Q (ram_74__7), .QB (\$dummy [1883]), .D (nx53200), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53201 (.Y (nx53200), .A0 (ram_74__7), .A1 (nx65476), .S0 (nx64026
             )) ;
    aoi22 ix62570 (.Y (nx62569), .A0 (ram_76__7), .A1 (nx64976), .B0 (ram_77__7)
          , .B1 (nx65014)) ;
    dffr reg_ram_76__7 (.Q (ram_76__7), .QB (\$dummy [1884]), .D (nx53180), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53181 (.Y (nx53180), .A0 (ram_76__7), .A1 (nx65476), .S0 (nx64018
             )) ;
    dffr reg_ram_77__7 (.Q (ram_77__7), .QB (\$dummy [1885]), .D (nx53170), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53171 (.Y (nx53170), .A0 (ram_77__7), .A1 (nx65476), .S0 (nx64014
             )) ;
    aoi22 ix62578 (.Y (nx62577), .A0 (ram_79__7), .A1 (nx65052), .B0 (ram_78__7)
          , .B1 (nx65090)) ;
    dffr reg_ram_79__7 (.Q (ram_79__7), .QB (\$dummy [1886]), .D (nx53150), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53151 (.Y (nx53150), .A0 (ram_79__7), .A1 (nx65476), .S0 (nx64006
             )) ;
    dffr reg_ram_78__7 (.Q (ram_78__7), .QB (\$dummy [1887]), .D (nx53160), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53161 (.Y (nx53160), .A0 (ram_78__7), .A1 (nx65476), .S0 (nx64010
             )) ;
    oai21 ix62586 (.Y (nx62585), .A0 (nx22156), .A1 (nx22078), .B0 (nx66144)) ;
    nand04 ix22157 (.Y (nx22156), .A0 (nx62588), .A1 (nx62596), .A2 (nx62604), .A3 (
           nx62612)) ;
    aoi22 ix62589 (.Y (nx62588), .A0 (ram_48__7), .A1 (nx64522), .B0 (ram_49__7)
          , .B1 (nx64560)) ;
    dffr reg_ram_48__7 (.Q (ram_48__7), .QB (\$dummy [1888]), .D (nx53140), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53141 (.Y (nx53140), .A0 (ram_48__7), .A1 (nx65476), .S0 (nx63996
             )) ;
    dffr reg_ram_49__7 (.Q (ram_49__7), .QB (\$dummy [1889]), .D (nx53130), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53131 (.Y (nx53130), .A0 (ram_49__7), .A1 (nx65476), .S0 (nx63992
             )) ;
    aoi22 ix62597 (.Y (nx62596), .A0 (ram_51__7), .A1 (nx64598), .B0 (ram_50__7)
          , .B1 (nx64636)) ;
    dffr reg_ram_51__7 (.Q (ram_51__7), .QB (\$dummy [1890]), .D (nx53110), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53111 (.Y (nx53110), .A0 (ram_51__7), .A1 (nx65478), .S0 (nx63984
             )) ;
    dffr reg_ram_50__7 (.Q (ram_50__7), .QB (\$dummy [1891]), .D (nx53120), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53121 (.Y (nx53120), .A0 (ram_50__7), .A1 (nx65478), .S0 (nx63988
             )) ;
    aoi22 ix62605 (.Y (nx62604), .A0 (ram_52__7), .A1 (nx64674), .B0 (ram_53__7)
          , .B1 (nx64712)) ;
    dffr reg_ram_52__7 (.Q (ram_52__7), .QB (\$dummy [1892]), .D (nx53100), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53101 (.Y (nx53100), .A0 (ram_52__7), .A1 (nx65478), .S0 (nx63980
             )) ;
    dffr reg_ram_53__7 (.Q (ram_53__7), .QB (\$dummy [1893]), .D (nx53090), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53091 (.Y (nx53090), .A0 (ram_53__7), .A1 (nx65478), .S0 (nx63976
             )) ;
    aoi22 ix62613 (.Y (nx62612), .A0 (ram_55__7), .A1 (nx64750), .B0 (ram_54__7)
          , .B1 (nx64788)) ;
    dffr reg_ram_55__7 (.Q (ram_55__7), .QB (\$dummy [1894]), .D (nx53070), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53071 (.Y (nx53070), .A0 (ram_55__7), .A1 (nx65478), .S0 (nx63968
             )) ;
    dffr reg_ram_54__7 (.Q (ram_54__7), .QB (\$dummy [1895]), .D (nx53080), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53081 (.Y (nx53080), .A0 (ram_54__7), .A1 (nx65478), .S0 (nx63972
             )) ;
    nand04 ix22079 (.Y (nx22078), .A0 (nx62621), .A1 (nx62629), .A2 (nx62637), .A3 (
           nx62645)) ;
    aoi22 ix62622 (.Y (nx62621), .A0 (ram_56__7), .A1 (nx64826), .B0 (ram_57__7)
          , .B1 (nx64864)) ;
    dffr reg_ram_56__7 (.Q (ram_56__7), .QB (\$dummy [1896]), .D (nx53060), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53061 (.Y (nx53060), .A0 (ram_56__7), .A1 (nx65478), .S0 (nx63964
             )) ;
    dffr reg_ram_57__7 (.Q (ram_57__7), .QB (\$dummy [1897]), .D (nx53050), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53051 (.Y (nx53050), .A0 (ram_57__7), .A1 (nx65480), .S0 (nx63960
             )) ;
    aoi22 ix62630 (.Y (nx62629), .A0 (ram_59__7), .A1 (nx64902), .B0 (ram_58__7)
          , .B1 (nx64940)) ;
    dffr reg_ram_59__7 (.Q (ram_59__7), .QB (\$dummy [1898]), .D (nx53030), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53031 (.Y (nx53030), .A0 (ram_59__7), .A1 (nx65480), .S0 (nx63952
             )) ;
    dffr reg_ram_58__7 (.Q (ram_58__7), .QB (\$dummy [1899]), .D (nx53040), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53041 (.Y (nx53040), .A0 (ram_58__7), .A1 (nx65480), .S0 (nx63956
             )) ;
    aoi22 ix62638 (.Y (nx62637), .A0 (ram_60__7), .A1 (nx64978), .B0 (ram_61__7)
          , .B1 (nx65016)) ;
    dffr reg_ram_60__7 (.Q (ram_60__7), .QB (\$dummy [1900]), .D (nx53020), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53021 (.Y (nx53020), .A0 (ram_60__7), .A1 (nx65480), .S0 (nx63948
             )) ;
    dffr reg_ram_61__7 (.Q (ram_61__7), .QB (\$dummy [1901]), .D (nx53010), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53011 (.Y (nx53010), .A0 (ram_61__7), .A1 (nx65480), .S0 (nx63944
             )) ;
    aoi22 ix62646 (.Y (nx62645), .A0 (ram_63__7), .A1 (nx65054), .B0 (ram_62__7)
          , .B1 (nx65092)) ;
    dffr reg_ram_63__7 (.Q (ram_63__7), .QB (\$dummy [1902]), .D (nx52990), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52991 (.Y (nx52990), .A0 (ram_63__7), .A1 (nx65480), .S0 (nx63936
             )) ;
    dffr reg_ram_62__7 (.Q (ram_62__7), .QB (\$dummy [1903]), .D (nx53000), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix53001 (.Y (nx53000), .A0 (ram_62__7), .A1 (nx65480), .S0 (nx63940
             )) ;
    oai21 ix62654 (.Y (nx62653), .A0 (nx21994), .A1 (nx21916), .B0 (nx66148)) ;
    nand04 ix21995 (.Y (nx21994), .A0 (nx62656), .A1 (nx62664), .A2 (nx62672), .A3 (
           nx62680)) ;
    aoi22 ix62657 (.Y (nx62656), .A0 (ram_32__7), .A1 (nx64522), .B0 (ram_33__7)
          , .B1 (nx64560)) ;
    dffr reg_ram_32__7 (.Q (ram_32__7), .QB (\$dummy [1904]), .D (nx52980), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52981 (.Y (nx52980), .A0 (ram_32__7), .A1 (nx65482), .S0 (nx63926
             )) ;
    dffr reg_ram_33__7 (.Q (ram_33__7), .QB (\$dummy [1905]), .D (nx52970), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52971 (.Y (nx52970), .A0 (ram_33__7), .A1 (nx65482), .S0 (nx63922
             )) ;
    aoi22 ix62665 (.Y (nx62664), .A0 (ram_35__7), .A1 (nx64598), .B0 (ram_34__7)
          , .B1 (nx64636)) ;
    dffr reg_ram_35__7 (.Q (ram_35__7), .QB (\$dummy [1906]), .D (nx52950), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52951 (.Y (nx52950), .A0 (ram_35__7), .A1 (nx65482), .S0 (nx63914
             )) ;
    dffr reg_ram_34__7 (.Q (ram_34__7), .QB (\$dummy [1907]), .D (nx52960), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52961 (.Y (nx52960), .A0 (ram_34__7), .A1 (nx65482), .S0 (nx63918
             )) ;
    aoi22 ix62673 (.Y (nx62672), .A0 (ram_36__7), .A1 (nx64674), .B0 (ram_37__7)
          , .B1 (nx64712)) ;
    dffr reg_ram_36__7 (.Q (ram_36__7), .QB (\$dummy [1908]), .D (nx52940), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52941 (.Y (nx52940), .A0 (ram_36__7), .A1 (nx65482), .S0 (nx63910
             )) ;
    dffr reg_ram_37__7 (.Q (ram_37__7), .QB (\$dummy [1909]), .D (nx52930), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52931 (.Y (nx52930), .A0 (ram_37__7), .A1 (nx65482), .S0 (nx63906
             )) ;
    aoi22 ix62681 (.Y (nx62680), .A0 (ram_39__7), .A1 (nx64750), .B0 (ram_38__7)
          , .B1 (nx64788)) ;
    dffr reg_ram_39__7 (.Q (ram_39__7), .QB (\$dummy [1910]), .D (nx52910), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52911 (.Y (nx52910), .A0 (ram_39__7), .A1 (nx65482), .S0 (nx63898
             )) ;
    dffr reg_ram_38__7 (.Q (ram_38__7), .QB (\$dummy [1911]), .D (nx52920), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52921 (.Y (nx52920), .A0 (ram_38__7), .A1 (nx65484), .S0 (nx63902
             )) ;
    nand04 ix21917 (.Y (nx21916), .A0 (nx62689), .A1 (nx62697), .A2 (nx62705), .A3 (
           nx62713)) ;
    aoi22 ix62690 (.Y (nx62689), .A0 (ram_40__7), .A1 (nx64826), .B0 (ram_41__7)
          , .B1 (nx64864)) ;
    dffr reg_ram_40__7 (.Q (ram_40__7), .QB (\$dummy [1912]), .D (nx52900), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52901 (.Y (nx52900), .A0 (ram_40__7), .A1 (nx65484), .S0 (nx63894
             )) ;
    dffr reg_ram_41__7 (.Q (ram_41__7), .QB (\$dummy [1913]), .D (nx52890), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52891 (.Y (nx52890), .A0 (ram_41__7), .A1 (nx65484), .S0 (nx63890
             )) ;
    aoi22 ix62698 (.Y (nx62697), .A0 (ram_43__7), .A1 (nx64902), .B0 (ram_42__7)
          , .B1 (nx64940)) ;
    dffr reg_ram_43__7 (.Q (ram_43__7), .QB (\$dummy [1914]), .D (nx52870), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52871 (.Y (nx52870), .A0 (ram_43__7), .A1 (nx65484), .S0 (nx63882
             )) ;
    dffr reg_ram_42__7 (.Q (ram_42__7), .QB (\$dummy [1915]), .D (nx52880), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52881 (.Y (nx52880), .A0 (ram_42__7), .A1 (nx65484), .S0 (nx63886
             )) ;
    aoi22 ix62706 (.Y (nx62705), .A0 (ram_44__7), .A1 (nx64978), .B0 (ram_45__7)
          , .B1 (nx65016)) ;
    dffr reg_ram_44__7 (.Q (ram_44__7), .QB (\$dummy [1916]), .D (nx52860), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52861 (.Y (nx52860), .A0 (ram_44__7), .A1 (nx65484), .S0 (nx63878
             )) ;
    dffr reg_ram_45__7 (.Q (ram_45__7), .QB (\$dummy [1917]), .D (nx52850), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52851 (.Y (nx52850), .A0 (ram_45__7), .A1 (nx65484), .S0 (nx63874
             )) ;
    aoi22 ix62714 (.Y (nx62713), .A0 (ram_47__7), .A1 (nx65054), .B0 (ram_46__7)
          , .B1 (nx65092)) ;
    dffr reg_ram_47__7 (.Q (ram_47__7), .QB (\$dummy [1918]), .D (nx52830), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52831 (.Y (nx52830), .A0 (ram_47__7), .A1 (nx65486), .S0 (nx63866
             )) ;
    dffr reg_ram_46__7 (.Q (ram_46__7), .QB (\$dummy [1919]), .D (nx52840), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52841 (.Y (nx52840), .A0 (ram_46__7), .A1 (nx65486), .S0 (nx63870
             )) ;
    nand04 ix21837 (.Y (nx21836), .A0 (nx62722), .A1 (nx62790), .A2 (nx62858), .A3 (
           nx62926)) ;
    oai21 ix62723 (.Y (nx62722), .A0 (nx21826), .A1 (nx21748), .B0 (nx66152)) ;
    nand04 ix21827 (.Y (nx21826), .A0 (nx62725), .A1 (nx62733), .A2 (nx62741), .A3 (
           nx62749)) ;
    aoi22 ix62726 (.Y (nx62725), .A0 (ram_16__7), .A1 (nx64522), .B0 (ram_17__7)
          , .B1 (nx64560)) ;
    dffr reg_ram_16__7 (.Q (ram_16__7), .QB (\$dummy [1920]), .D (nx52820), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52821 (.Y (nx52820), .A0 (ram_16__7), .A1 (nx65486), .S0 (nx63856
             )) ;
    dffr reg_ram_17__7 (.Q (ram_17__7), .QB (\$dummy [1921]), .D (nx52810), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52811 (.Y (nx52810), .A0 (ram_17__7), .A1 (nx65486), .S0 (nx63852
             )) ;
    aoi22 ix62734 (.Y (nx62733), .A0 (ram_19__7), .A1 (nx64598), .B0 (ram_18__7)
          , .B1 (nx64636)) ;
    dffr reg_ram_19__7 (.Q (ram_19__7), .QB (\$dummy [1922]), .D (nx52790), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52791 (.Y (nx52790), .A0 (ram_19__7), .A1 (nx65486), .S0 (nx63844
             )) ;
    dffr reg_ram_18__7 (.Q (ram_18__7), .QB (\$dummy [1923]), .D (nx52800), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52801 (.Y (nx52800), .A0 (ram_18__7), .A1 (nx65486), .S0 (nx63848
             )) ;
    aoi22 ix62742 (.Y (nx62741), .A0 (ram_20__7), .A1 (nx64674), .B0 (ram_21__7)
          , .B1 (nx64712)) ;
    dffr reg_ram_20__7 (.Q (ram_20__7), .QB (\$dummy [1924]), .D (nx52780), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52781 (.Y (nx52780), .A0 (ram_20__7), .A1 (nx65486), .S0 (nx63840
             )) ;
    dffr reg_ram_21__7 (.Q (ram_21__7), .QB (\$dummy [1925]), .D (nx52770), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52771 (.Y (nx52770), .A0 (ram_21__7), .A1 (nx65488), .S0 (nx63836
             )) ;
    aoi22 ix62750 (.Y (nx62749), .A0 (ram_23__7), .A1 (nx64750), .B0 (ram_22__7)
          , .B1 (nx64788)) ;
    dffr reg_ram_23__7 (.Q (ram_23__7), .QB (\$dummy [1926]), .D (nx52750), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52751 (.Y (nx52750), .A0 (ram_23__7), .A1 (nx65488), .S0 (nx63828
             )) ;
    dffr reg_ram_22__7 (.Q (ram_22__7), .QB (\$dummy [1927]), .D (nx52760), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52761 (.Y (nx52760), .A0 (ram_22__7), .A1 (nx65488), .S0 (nx63832
             )) ;
    nand04 ix21749 (.Y (nx21748), .A0 (nx62758), .A1 (nx62766), .A2 (nx62774), .A3 (
           nx62782)) ;
    aoi22 ix62759 (.Y (nx62758), .A0 (ram_24__7), .A1 (nx64826), .B0 (ram_25__7)
          , .B1 (nx64864)) ;
    dffr reg_ram_24__7 (.Q (ram_24__7), .QB (\$dummy [1928]), .D (nx52740), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52741 (.Y (nx52740), .A0 (ram_24__7), .A1 (nx65488), .S0 (nx63824
             )) ;
    dffr reg_ram_25__7 (.Q (ram_25__7), .QB (\$dummy [1929]), .D (nx52730), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52731 (.Y (nx52730), .A0 (ram_25__7), .A1 (nx65488), .S0 (nx63820
             )) ;
    aoi22 ix62767 (.Y (nx62766), .A0 (ram_27__7), .A1 (nx64902), .B0 (ram_26__7)
          , .B1 (nx64940)) ;
    dffr reg_ram_27__7 (.Q (ram_27__7), .QB (\$dummy [1930]), .D (nx52710), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52711 (.Y (nx52710), .A0 (ram_27__7), .A1 (nx65488), .S0 (nx63812
             )) ;
    dffr reg_ram_26__7 (.Q (ram_26__7), .QB (\$dummy [1931]), .D (nx52720), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52721 (.Y (nx52720), .A0 (ram_26__7), .A1 (nx65488), .S0 (nx63816
             )) ;
    aoi22 ix62775 (.Y (nx62774), .A0 (ram_28__7), .A1 (nx64978), .B0 (ram_29__7)
          , .B1 (nx65016)) ;
    dffr reg_ram_28__7 (.Q (ram_28__7), .QB (\$dummy [1932]), .D (nx52700), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52701 (.Y (nx52700), .A0 (ram_28__7), .A1 (nx65490), .S0 (nx63808
             )) ;
    dffr reg_ram_29__7 (.Q (ram_29__7), .QB (\$dummy [1933]), .D (nx52690), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52691 (.Y (nx52690), .A0 (ram_29__7), .A1 (nx65490), .S0 (nx63804
             )) ;
    aoi22 ix62783 (.Y (nx62782), .A0 (ram_31__7), .A1 (nx65054), .B0 (ram_30__7)
          , .B1 (nx65092)) ;
    dffr reg_ram_31__7 (.Q (ram_31__7), .QB (\$dummy [1934]), .D (nx52670), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52671 (.Y (nx52670), .A0 (ram_31__7), .A1 (nx65490), .S0 (nx63796
             )) ;
    dffr reg_ram_30__7 (.Q (ram_30__7), .QB (\$dummy [1935]), .D (nx52680), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52681 (.Y (nx52680), .A0 (ram_30__7), .A1 (nx65490), .S0 (nx63800
             )) ;
    oai21 ix62791 (.Y (nx62790), .A0 (nx21664), .A1 (nx21586), .B0 (nx65144)) ;
    nand04 ix21665 (.Y (nx21664), .A0 (nx62793), .A1 (nx62801), .A2 (nx62809), .A3 (
           nx62817)) ;
    aoi22 ix62794 (.Y (nx62793), .A0 (ram_0__7), .A1 (nx64522), .B0 (ram_1__7), 
          .B1 (nx64560)) ;
    dffr reg_ram_0__7 (.Q (ram_0__7), .QB (\$dummy [1936]), .D (nx52660), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52661 (.Y (nx52660), .A0 (nx65490), .A1 (ram_0__7), .S0 (nx65134)
             ) ;
    dffr reg_ram_1__7 (.Q (ram_1__7), .QB (\$dummy [1937]), .D (nx52650), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52651 (.Y (nx52650), .A0 (nx65490), .A1 (ram_1__7), .S0 (nx65148)
             ) ;
    aoi22 ix62802 (.Y (nx62801), .A0 (ram_3__7), .A1 (nx64598), .B0 (ram_2__7), 
          .B1 (nx64636)) ;
    dffr reg_ram_3__7 (.Q (ram_3__7), .QB (\$dummy [1938]), .D (nx52630), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52631 (.Y (nx52630), .A0 (nx65490), .A1 (ram_3__7), .S0 (nx65152)
             ) ;
    dffr reg_ram_2__7 (.Q (ram_2__7), .QB (\$dummy [1939]), .D (nx52640), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52641 (.Y (nx52640), .A0 (nx65492), .A1 (ram_2__7), .S0 (nx65156)
             ) ;
    aoi22 ix62810 (.Y (nx62809), .A0 (ram_4__7), .A1 (nx64674), .B0 (ram_5__7), 
          .B1 (nx64712)) ;
    dffr reg_ram_4__7 (.Q (ram_4__7), .QB (\$dummy [1940]), .D (nx52620), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52621 (.Y (nx52620), .A0 (nx65492), .A1 (ram_4__7), .S0 (nx65160)
             ) ;
    dffr reg_ram_5__7 (.Q (ram_5__7), .QB (\$dummy [1941]), .D (nx52610), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52611 (.Y (nx52610), .A0 (nx65492), .A1 (ram_5__7), .S0 (nx65164)
             ) ;
    aoi22 ix62818 (.Y (nx62817), .A0 (ram_7__7), .A1 (nx64750), .B0 (ram_6__7), 
          .B1 (nx64788)) ;
    dffr reg_ram_7__7 (.Q (ram_7__7), .QB (\$dummy [1942]), .D (nx52590), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52591 (.Y (nx52590), .A0 (nx65492), .A1 (ram_7__7), .S0 (nx65168)
             ) ;
    dffr reg_ram_6__7 (.Q (ram_6__7), .QB (\$dummy [1943]), .D (nx52600), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52601 (.Y (nx52600), .A0 (nx65492), .A1 (ram_6__7), .S0 (nx65172)
             ) ;
    nand04 ix21587 (.Y (nx21586), .A0 (nx62826), .A1 (nx62834), .A2 (nx62842), .A3 (
           nx62850)) ;
    aoi22 ix62827 (.Y (nx62826), .A0 (ram_8__7), .A1 (nx64826), .B0 (ram_9__7), 
          .B1 (nx64864)) ;
    dffr reg_ram_8__7 (.Q (ram_8__7), .QB (\$dummy [1944]), .D (nx52580), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52581 (.Y (nx52580), .A0 (nx65492), .A1 (ram_8__7), .S0 (nx65176)
             ) ;
    dffr reg_ram_9__7 (.Q (ram_9__7), .QB (\$dummy [1945]), .D (nx52570), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52571 (.Y (nx52570), .A0 (nx65492), .A1 (ram_9__7), .S0 (nx65180)
             ) ;
    aoi22 ix62835 (.Y (nx62834), .A0 (ram_11__7), .A1 (nx64902), .B0 (ram_10__7)
          , .B1 (nx64940)) ;
    dffr reg_ram_11__7 (.Q (ram_11__7), .QB (\$dummy [1946]), .D (nx52550), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52551 (.Y (nx52550), .A0 (nx65494), .A1 (ram_11__7), .S0 (nx65184
             )) ;
    dffr reg_ram_10__7 (.Q (ram_10__7), .QB (\$dummy [1947]), .D (nx52560), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52561 (.Y (nx52560), .A0 (nx65494), .A1 (ram_10__7), .S0 (nx65188
             )) ;
    aoi22 ix62843 (.Y (nx62842), .A0 (ram_12__7), .A1 (nx64978), .B0 (ram_13__7)
          , .B1 (nx65016)) ;
    dffr reg_ram_12__7 (.Q (ram_12__7), .QB (\$dummy [1948]), .D (nx52540), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52541 (.Y (nx52540), .A0 (nx65494), .A1 (ram_12__7), .S0 (nx65192
             )) ;
    dffr reg_ram_13__7 (.Q (ram_13__7), .QB (\$dummy [1949]), .D (nx52530), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52531 (.Y (nx52530), .A0 (nx65494), .A1 (ram_13__7), .S0 (nx65196
             )) ;
    aoi22 ix62851 (.Y (nx62850), .A0 (ram_15__7), .A1 (nx65054), .B0 (ram_14__7)
          , .B1 (nx65092)) ;
    dffr reg_ram_15__7 (.Q (ram_15__7), .QB (\$dummy [1950]), .D (nx52510), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52511 (.Y (nx52510), .A0 (nx65494), .A1 (ram_15__7), .S0 (nx65200
             )) ;
    dffr reg_ram_14__7 (.Q (ram_14__7), .QB (\$dummy [1951]), .D (nx52520), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52521 (.Y (nx52520), .A0 (nx65494), .A1 (ram_14__7), .S0 (nx65204
             )) ;
    oai21 ix62859 (.Y (nx62858), .A0 (nx21500), .A1 (nx21422), .B0 (nx66156)) ;
    nand04 ix21501 (.Y (nx21500), .A0 (nx62861), .A1 (nx62869), .A2 (nx62877), .A3 (
           nx62885)) ;
    aoi22 ix62862 (.Y (nx62861), .A0 (ram_96__7), .A1 (nx64522), .B0 (ram_97__7)
          , .B1 (nx64560)) ;
    dffr reg_ram_96__7 (.Q (ram_96__7), .QB (\$dummy [1952]), .D (nx52500), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52501 (.Y (nx52500), .A0 (ram_96__7), .A1 (nx65494), .S0 (nx63786
             )) ;
    dffr reg_ram_97__7 (.Q (ram_97__7), .QB (\$dummy [1953]), .D (nx52490), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52491 (.Y (nx52490), .A0 (ram_97__7), .A1 (nx65496), .S0 (nx63782
             )) ;
    aoi22 ix62870 (.Y (nx62869), .A0 (ram_99__7), .A1 (nx64598), .B0 (ram_98__7)
          , .B1 (nx64636)) ;
    dffr reg_ram_99__7 (.Q (ram_99__7), .QB (\$dummy [1954]), .D (nx52470), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52471 (.Y (nx52470), .A0 (ram_99__7), .A1 (nx65496), .S0 (nx63774
             )) ;
    dffr reg_ram_98__7 (.Q (ram_98__7), .QB (\$dummy [1955]), .D (nx52480), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52481 (.Y (nx52480), .A0 (ram_98__7), .A1 (nx65496), .S0 (nx63778
             )) ;
    aoi22 ix62878 (.Y (nx62877), .A0 (ram_100__7), .A1 (nx64674), .B0 (
          ram_101__7), .B1 (nx64712)) ;
    dffr reg_ram_100__7 (.Q (ram_100__7), .QB (\$dummy [1956]), .D (nx52460), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52461 (.Y (nx52460), .A0 (ram_100__7), .A1 (nx65496), .S0 (
             nx63770)) ;
    dffr reg_ram_101__7 (.Q (ram_101__7), .QB (\$dummy [1957]), .D (nx52450), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52451 (.Y (nx52450), .A0 (ram_101__7), .A1 (nx65496), .S0 (
             nx63766)) ;
    aoi22 ix62886 (.Y (nx62885), .A0 (ram_103__7), .A1 (nx64750), .B0 (
          ram_102__7), .B1 (nx64788)) ;
    dffr reg_ram_103__7 (.Q (ram_103__7), .QB (\$dummy [1958]), .D (nx52430), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52431 (.Y (nx52430), .A0 (ram_103__7), .A1 (nx65496), .S0 (
             nx63758)) ;
    dffr reg_ram_102__7 (.Q (ram_102__7), .QB (\$dummy [1959]), .D (nx52440), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52441 (.Y (nx52440), .A0 (ram_102__7), .A1 (nx65496), .S0 (
             nx63762)) ;
    nand04 ix21423 (.Y (nx21422), .A0 (nx62894), .A1 (nx62902), .A2 (nx62910), .A3 (
           nx62918)) ;
    aoi22 ix62895 (.Y (nx62894), .A0 (ram_104__7), .A1 (nx64826), .B0 (
          ram_105__7), .B1 (nx64864)) ;
    dffr reg_ram_104__7 (.Q (ram_104__7), .QB (\$dummy [1960]), .D (nx52420), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52421 (.Y (nx52420), .A0 (ram_104__7), .A1 (nx65498), .S0 (
             nx63754)) ;
    dffr reg_ram_105__7 (.Q (ram_105__7), .QB (\$dummy [1961]), .D (nx52410), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52411 (.Y (nx52410), .A0 (ram_105__7), .A1 (nx65498), .S0 (
             nx63750)) ;
    aoi22 ix62903 (.Y (nx62902), .A0 (ram_107__7), .A1 (nx64902), .B0 (
          ram_106__7), .B1 (nx64940)) ;
    dffr reg_ram_107__7 (.Q (ram_107__7), .QB (\$dummy [1962]), .D (nx52390), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52391 (.Y (nx52390), .A0 (ram_107__7), .A1 (nx65498), .S0 (
             nx63742)) ;
    dffr reg_ram_106__7 (.Q (ram_106__7), .QB (\$dummy [1963]), .D (nx52400), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52401 (.Y (nx52400), .A0 (ram_106__7), .A1 (nx65498), .S0 (
             nx63746)) ;
    aoi22 ix62911 (.Y (nx62910), .A0 (ram_108__7), .A1 (nx64978), .B0 (
          ram_109__7), .B1 (nx65016)) ;
    dffr reg_ram_108__7 (.Q (ram_108__7), .QB (\$dummy [1964]), .D (nx52380), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52381 (.Y (nx52380), .A0 (ram_108__7), .A1 (nx65498), .S0 (
             nx63738)) ;
    dffr reg_ram_109__7 (.Q (ram_109__7), .QB (\$dummy [1965]), .D (nx52370), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52371 (.Y (nx52370), .A0 (ram_109__7), .A1 (nx65498), .S0 (
             nx63734)) ;
    aoi22 ix62919 (.Y (nx62918), .A0 (ram_111__7), .A1 (nx65054), .B0 (
          ram_110__7), .B1 (nx65092)) ;
    dffr reg_ram_111__7 (.Q (ram_111__7), .QB (\$dummy [1966]), .D (nx52350), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52351 (.Y (nx52350), .A0 (ram_111__7), .A1 (nx65498), .S0 (
             nx63726)) ;
    dffr reg_ram_110__7 (.Q (ram_110__7), .QB (\$dummy [1967]), .D (nx52360), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52361 (.Y (nx52360), .A0 (ram_110__7), .A1 (nx65500), .S0 (
             nx63730)) ;
    oai21 ix62927 (.Y (nx62926), .A0 (nx21338), .A1 (nx21260), .B0 (nx66160)) ;
    nand04 ix21339 (.Y (nx21338), .A0 (nx62929), .A1 (nx62937), .A2 (nx62945), .A3 (
           nx62953)) ;
    aoi22 ix62930 (.Y (nx62929), .A0 (ram_112__7), .A1 (nx64522), .B0 (
          ram_113__7), .B1 (nx64560)) ;
    dffr reg_ram_112__7 (.Q (ram_112__7), .QB (\$dummy [1968]), .D (nx52340), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52341 (.Y (nx52340), .A0 (ram_112__7), .A1 (nx65500), .S0 (
             nx63716)) ;
    dffr reg_ram_113__7 (.Q (ram_113__7), .QB (\$dummy [1969]), .D (nx52330), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52331 (.Y (nx52330), .A0 (ram_113__7), .A1 (nx65500), .S0 (
             nx63712)) ;
    aoi22 ix62938 (.Y (nx62937), .A0 (ram_115__7), .A1 (nx64598), .B0 (
          ram_114__7), .B1 (nx64636)) ;
    dffr reg_ram_115__7 (.Q (ram_115__7), .QB (\$dummy [1970]), .D (nx52310), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52311 (.Y (nx52310), .A0 (ram_115__7), .A1 (nx65500), .S0 (
             nx63704)) ;
    dffr reg_ram_114__7 (.Q (ram_114__7), .QB (\$dummy [1971]), .D (nx52320), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52321 (.Y (nx52320), .A0 (ram_114__7), .A1 (nx65500), .S0 (
             nx63708)) ;
    aoi22 ix62946 (.Y (nx62945), .A0 (ram_116__7), .A1 (nx64674), .B0 (
          ram_117__7), .B1 (nx64712)) ;
    dffr reg_ram_116__7 (.Q (ram_116__7), .QB (\$dummy [1972]), .D (nx52300), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52301 (.Y (nx52300), .A0 (ram_116__7), .A1 (nx65500), .S0 (
             nx63700)) ;
    dffr reg_ram_117__7 (.Q (ram_117__7), .QB (\$dummy [1973]), .D (nx52290), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52291 (.Y (nx52290), .A0 (ram_117__7), .A1 (nx65500), .S0 (
             nx63696)) ;
    aoi22 ix62954 (.Y (nx62953), .A0 (ram_119__7), .A1 (nx64750), .B0 (
          ram_118__7), .B1 (nx64788)) ;
    dffr reg_ram_119__7 (.Q (ram_119__7), .QB (\$dummy [1974]), .D (nx52270), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52271 (.Y (nx52270), .A0 (ram_119__7), .A1 (nx65502), .S0 (
             nx63688)) ;
    dffr reg_ram_118__7 (.Q (ram_118__7), .QB (\$dummy [1975]), .D (nx52280), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52281 (.Y (nx52280), .A0 (ram_118__7), .A1 (nx65502), .S0 (
             nx63692)) ;
    nand04 ix21261 (.Y (nx21260), .A0 (nx62962), .A1 (nx62970), .A2 (nx62978), .A3 (
           nx62986)) ;
    aoi22 ix62963 (.Y (nx62962), .A0 (ram_120__7), .A1 (nx64826), .B0 (
          ram_121__7), .B1 (nx64864)) ;
    dffr reg_ram_120__7 (.Q (ram_120__7), .QB (\$dummy [1976]), .D (nx52260), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52261 (.Y (nx52260), .A0 (ram_120__7), .A1 (nx65502), .S0 (
             nx63684)) ;
    dffr reg_ram_121__7 (.Q (ram_121__7), .QB (\$dummy [1977]), .D (nx52250), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52251 (.Y (nx52250), .A0 (ram_121__7), .A1 (nx65502), .S0 (
             nx63680)) ;
    aoi22 ix62971 (.Y (nx62970), .A0 (ram_123__7), .A1 (nx64902), .B0 (
          ram_122__7), .B1 (nx64940)) ;
    dffr reg_ram_123__7 (.Q (ram_123__7), .QB (\$dummy [1978]), .D (nx52230), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52231 (.Y (nx52230), .A0 (ram_123__7), .A1 (nx65502), .S0 (
             nx63672)) ;
    dffr reg_ram_122__7 (.Q (ram_122__7), .QB (\$dummy [1979]), .D (nx52240), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52241 (.Y (nx52240), .A0 (ram_122__7), .A1 (nx65502), .S0 (
             nx63676)) ;
    aoi22 ix62979 (.Y (nx62978), .A0 (ram_124__7), .A1 (nx64978), .B0 (
          ram_125__7), .B1 (nx65016)) ;
    dffr reg_ram_124__7 (.Q (ram_124__7), .QB (\$dummy [1980]), .D (nx52220), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52221 (.Y (nx52220), .A0 (ram_124__7), .A1 (nx65502), .S0 (
             nx63668)) ;
    dffr reg_ram_125__7 (.Q (ram_125__7), .QB (\$dummy [1981]), .D (nx52210), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52211 (.Y (nx52210), .A0 (ram_125__7), .A1 (nx65504), .S0 (
             nx63664)) ;
    aoi22 ix62987 (.Y (nx62986), .A0 (ram_127__7), .A1 (nx65054), .B0 (
          ram_126__7), .B1 (nx65092)) ;
    dffr reg_ram_127__7 (.Q (ram_127__7), .QB (\$dummy [1982]), .D (nx52190), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52191 (.Y (nx52190), .A0 (ram_127__7), .A1 (nx65504), .S0 (
             nx63656)) ;
    dffr reg_ram_126__7 (.Q (ram_126__7), .QB (\$dummy [1983]), .D (nx52200), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52201 (.Y (nx52200), .A0 (ram_126__7), .A1 (nx65504), .S0 (
             nx63660)) ;
    nand04 ix21183 (.Y (nx21182), .A0 (nx62995), .A1 (nx63063), .A2 (nx63131), .A3 (
           nx63199)) ;
    oai21 ix62996 (.Y (nx62995), .A0 (nx21172), .A1 (nx21094), .B0 (nx66164)) ;
    nand04 ix21173 (.Y (nx21172), .A0 (nx62998), .A1 (nx63006), .A2 (nx63014), .A3 (
           nx63022)) ;
    aoi22 ix62999 (.Y (nx62998), .A0 (ram_128__7), .A1 (nx64522), .B0 (
          ram_129__7), .B1 (nx64560)) ;
    dffr reg_ram_128__7 (.Q (ram_128__7), .QB (\$dummy [1984]), .D (nx52180), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52181 (.Y (nx52180), .A0 (ram_128__7), .A1 (nx65504), .S0 (
             nx63646)) ;
    dffr reg_ram_129__7 (.Q (ram_129__7), .QB (\$dummy [1985]), .D (nx52170), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52171 (.Y (nx52170), .A0 (ram_129__7), .A1 (nx65504), .S0 (
             nx63642)) ;
    aoi22 ix63007 (.Y (nx63006), .A0 (ram_131__7), .A1 (nx64598), .B0 (
          ram_130__7), .B1 (nx64636)) ;
    dffr reg_ram_131__7 (.Q (ram_131__7), .QB (\$dummy [1986]), .D (nx52150), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52151 (.Y (nx52150), .A0 (ram_131__7), .A1 (nx65504), .S0 (
             nx63634)) ;
    dffr reg_ram_130__7 (.Q (ram_130__7), .QB (\$dummy [1987]), .D (nx52160), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52161 (.Y (nx52160), .A0 (ram_130__7), .A1 (nx65504), .S0 (
             nx63638)) ;
    aoi22 ix63015 (.Y (nx63014), .A0 (ram_132__7), .A1 (nx64674), .B0 (
          ram_133__7), .B1 (nx64712)) ;
    dffr reg_ram_132__7 (.Q (ram_132__7), .QB (\$dummy [1988]), .D (nx52140), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52141 (.Y (nx52140), .A0 (ram_132__7), .A1 (nx65506), .S0 (
             nx63630)) ;
    dffr reg_ram_133__7 (.Q (ram_133__7), .QB (\$dummy [1989]), .D (nx52130), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52131 (.Y (nx52130), .A0 (ram_133__7), .A1 (nx65506), .S0 (
             nx63626)) ;
    aoi22 ix63023 (.Y (nx63022), .A0 (ram_135__7), .A1 (nx64750), .B0 (
          ram_134__7), .B1 (nx64788)) ;
    dffr reg_ram_135__7 (.Q (ram_135__7), .QB (\$dummy [1990]), .D (nx52110), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52111 (.Y (nx52110), .A0 (ram_135__7), .A1 (nx65506), .S0 (
             nx63618)) ;
    dffr reg_ram_134__7 (.Q (ram_134__7), .QB (\$dummy [1991]), .D (nx52120), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52121 (.Y (nx52120), .A0 (ram_134__7), .A1 (nx65506), .S0 (
             nx63622)) ;
    nand04 ix21095 (.Y (nx21094), .A0 (nx63031), .A1 (nx63039), .A2 (nx63047), .A3 (
           nx63055)) ;
    aoi22 ix63032 (.Y (nx63031), .A0 (ram_136__7), .A1 (nx64826), .B0 (
          ram_137__7), .B1 (nx64864)) ;
    dffr reg_ram_136__7 (.Q (ram_136__7), .QB (\$dummy [1992]), .D (nx52100), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52101 (.Y (nx52100), .A0 (ram_136__7), .A1 (nx65506), .S0 (
             nx63614)) ;
    dffr reg_ram_137__7 (.Q (ram_137__7), .QB (\$dummy [1993]), .D (nx52090), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52091 (.Y (nx52090), .A0 (ram_137__7), .A1 (nx65506), .S0 (
             nx63610)) ;
    aoi22 ix63040 (.Y (nx63039), .A0 (ram_139__7), .A1 (nx64902), .B0 (
          ram_138__7), .B1 (nx64940)) ;
    dffr reg_ram_139__7 (.Q (ram_139__7), .QB (\$dummy [1994]), .D (nx52070), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52071 (.Y (nx52070), .A0 (ram_139__7), .A1 (nx65506), .S0 (
             nx63602)) ;
    dffr reg_ram_138__7 (.Q (ram_138__7), .QB (\$dummy [1995]), .D (nx52080), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52081 (.Y (nx52080), .A0 (ram_138__7), .A1 (nx65508), .S0 (
             nx63606)) ;
    aoi22 ix63048 (.Y (nx63047), .A0 (ram_140__7), .A1 (nx64978), .B0 (
          ram_141__7), .B1 (nx65016)) ;
    dffr reg_ram_140__7 (.Q (ram_140__7), .QB (\$dummy [1996]), .D (nx52060), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52061 (.Y (nx52060), .A0 (ram_140__7), .A1 (nx65508), .S0 (
             nx63598)) ;
    dffr reg_ram_141__7 (.Q (ram_141__7), .QB (\$dummy [1997]), .D (nx52050), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52051 (.Y (nx52050), .A0 (ram_141__7), .A1 (nx65508), .S0 (
             nx63594)) ;
    aoi22 ix63056 (.Y (nx63055), .A0 (ram_143__7), .A1 (nx65054), .B0 (
          ram_142__7), .B1 (nx65092)) ;
    dffr reg_ram_143__7 (.Q (ram_143__7), .QB (\$dummy [1998]), .D (nx52030), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52031 (.Y (nx52030), .A0 (ram_143__7), .A1 (nx65508), .S0 (
             nx63586)) ;
    dffr reg_ram_142__7 (.Q (ram_142__7), .QB (\$dummy [1999]), .D (nx52040), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52041 (.Y (nx52040), .A0 (ram_142__7), .A1 (nx65508), .S0 (
             nx63590)) ;
    oai21 ix63064 (.Y (nx63063), .A0 (nx21010), .A1 (nx20932), .B0 (nx66168)) ;
    nand04 ix21011 (.Y (nx21010), .A0 (nx63066), .A1 (nx63074), .A2 (nx63082), .A3 (
           nx63090)) ;
    aoi22 ix63067 (.Y (nx63066), .A0 (ram_144__7), .A1 (nx66056), .B0 (
          ram_145__7), .B1 (nx66060)) ;
    dffr reg_ram_144__7 (.Q (ram_144__7), .QB (\$dummy [2000]), .D (nx52020), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52021 (.Y (nx52020), .A0 (ram_144__7), .A1 (nx65508), .S0 (
             nx63576)) ;
    dffr reg_ram_145__7 (.Q (ram_145__7), .QB (\$dummy [2001]), .D (nx52010), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52011 (.Y (nx52010), .A0 (ram_145__7), .A1 (nx65508), .S0 (
             nx63572)) ;
    aoi22 ix63075 (.Y (nx63074), .A0 (ram_147__7), .A1 (nx66064), .B0 (
          ram_146__7), .B1 (nx66068)) ;
    dffr reg_ram_147__7 (.Q (ram_147__7), .QB (\$dummy [2002]), .D (nx51990), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51991 (.Y (nx51990), .A0 (ram_147__7), .A1 (nx65510), .S0 (
             nx63564)) ;
    dffr reg_ram_146__7 (.Q (ram_146__7), .QB (\$dummy [2003]), .D (nx52000), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix52001 (.Y (nx52000), .A0 (ram_146__7), .A1 (nx65510), .S0 (
             nx63568)) ;
    aoi22 ix63083 (.Y (nx63082), .A0 (ram_148__7), .A1 (nx66072), .B0 (
          ram_149__7), .B1 (nx66076)) ;
    dffr reg_ram_148__7 (.Q (ram_148__7), .QB (\$dummy [2004]), .D (nx51980), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51981 (.Y (nx51980), .A0 (ram_148__7), .A1 (nx65510), .S0 (
             nx63560)) ;
    dffr reg_ram_149__7 (.Q (ram_149__7), .QB (\$dummy [2005]), .D (nx51970), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51971 (.Y (nx51970), .A0 (ram_149__7), .A1 (nx65510), .S0 (
             nx63556)) ;
    aoi22 ix63091 (.Y (nx63090), .A0 (ram_151__7), .A1 (nx66080), .B0 (
          ram_150__7), .B1 (nx66084)) ;
    dffr reg_ram_151__7 (.Q (ram_151__7), .QB (\$dummy [2006]), .D (nx51950), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51951 (.Y (nx51950), .A0 (ram_151__7), .A1 (nx65510), .S0 (
             nx63548)) ;
    dffr reg_ram_150__7 (.Q (ram_150__7), .QB (\$dummy [2007]), .D (nx51960), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51961 (.Y (nx51960), .A0 (ram_150__7), .A1 (nx65510), .S0 (
             nx63552)) ;
    nand04 ix20933 (.Y (nx20932), .A0 (nx63099), .A1 (nx63107), .A2 (nx63115), .A3 (
           nx63123)) ;
    aoi22 ix63100 (.Y (nx63099), .A0 (ram_152__7), .A1 (nx66088), .B0 (
          ram_153__7), .B1 (nx66092)) ;
    dffr reg_ram_152__7 (.Q (ram_152__7), .QB (\$dummy [2008]), .D (nx51940), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51941 (.Y (nx51940), .A0 (ram_152__7), .A1 (nx65510), .S0 (
             nx63544)) ;
    dffr reg_ram_153__7 (.Q (ram_153__7), .QB (\$dummy [2009]), .D (nx51930), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51931 (.Y (nx51930), .A0 (ram_153__7), .A1 (nx65512), .S0 (
             nx63540)) ;
    aoi22 ix63108 (.Y (nx63107), .A0 (ram_155__7), .A1 (nx66096), .B0 (
          ram_154__7), .B1 (nx66100)) ;
    dffr reg_ram_155__7 (.Q (ram_155__7), .QB (\$dummy [2010]), .D (nx51910), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51911 (.Y (nx51910), .A0 (ram_155__7), .A1 (nx65512), .S0 (
             nx63532)) ;
    dffr reg_ram_154__7 (.Q (ram_154__7), .QB (\$dummy [2011]), .D (nx51920), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51921 (.Y (nx51920), .A0 (ram_154__7), .A1 (nx65512), .S0 (
             nx63536)) ;
    aoi22 ix63116 (.Y (nx63115), .A0 (ram_156__7), .A1 (nx66104), .B0 (
          ram_157__7), .B1 (nx66108)) ;
    dffr reg_ram_156__7 (.Q (ram_156__7), .QB (\$dummy [2012]), .D (nx51900), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51901 (.Y (nx51900), .A0 (ram_156__7), .A1 (nx65512), .S0 (
             nx63528)) ;
    dffr reg_ram_157__7 (.Q (ram_157__7), .QB (\$dummy [2013]), .D (nx51890), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51891 (.Y (nx51890), .A0 (ram_157__7), .A1 (nx65512), .S0 (
             nx63524)) ;
    aoi22 ix63124 (.Y (nx63123), .A0 (ram_159__7), .A1 (nx66112), .B0 (
          ram_158__7), .B1 (nx66116)) ;
    dffr reg_ram_159__7 (.Q (ram_159__7), .QB (\$dummy [2014]), .D (nx51870), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51871 (.Y (nx51870), .A0 (ram_159__7), .A1 (nx65512), .S0 (
             nx63516)) ;
    dffr reg_ram_158__7 (.Q (ram_158__7), .QB (\$dummy [2015]), .D (nx51880), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51881 (.Y (nx51880), .A0 (ram_158__7), .A1 (nx65512), .S0 (
             nx63520)) ;
    oai21 ix63132 (.Y (nx63131), .A0 (nx20846), .A1 (nx20768), .B0 (nx66172)) ;
    nand04 ix20847 (.Y (nx20846), .A0 (nx63134), .A1 (nx63142), .A2 (nx63150), .A3 (
           nx63158)) ;
    aoi22 ix63135 (.Y (nx63134), .A0 (ram_160__7), .A1 (nx66056), .B0 (
          ram_161__7), .B1 (nx66060)) ;
    dffr reg_ram_160__7 (.Q (ram_160__7), .QB (\$dummy [2016]), .D (nx51860), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51861 (.Y (nx51860), .A0 (ram_160__7), .A1 (nx65514), .S0 (
             nx63506)) ;
    dffr reg_ram_161__7 (.Q (ram_161__7), .QB (\$dummy [2017]), .D (nx51850), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51851 (.Y (nx51850), .A0 (ram_161__7), .A1 (nx65514), .S0 (
             nx63502)) ;
    aoi22 ix63143 (.Y (nx63142), .A0 (ram_163__7), .A1 (nx66064), .B0 (
          ram_162__7), .B1 (nx66068)) ;
    dffr reg_ram_163__7 (.Q (ram_163__7), .QB (\$dummy [2018]), .D (nx51830), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51831 (.Y (nx51830), .A0 (ram_163__7), .A1 (nx65514), .S0 (
             nx63494)) ;
    dffr reg_ram_162__7 (.Q (ram_162__7), .QB (\$dummy [2019]), .D (nx51840), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51841 (.Y (nx51840), .A0 (ram_162__7), .A1 (nx65514), .S0 (
             nx63498)) ;
    aoi22 ix63151 (.Y (nx63150), .A0 (ram_164__7), .A1 (nx66072), .B0 (
          ram_165__7), .B1 (nx66076)) ;
    dffr reg_ram_164__7 (.Q (ram_164__7), .QB (\$dummy [2020]), .D (nx51820), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51821 (.Y (nx51820), .A0 (ram_164__7), .A1 (nx65514), .S0 (
             nx63490)) ;
    dffr reg_ram_165__7 (.Q (ram_165__7), .QB (\$dummy [2021]), .D (nx51810), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51811 (.Y (nx51810), .A0 (ram_165__7), .A1 (nx65514), .S0 (
             nx63486)) ;
    aoi22 ix63159 (.Y (nx63158), .A0 (ram_167__7), .A1 (nx66080), .B0 (
          ram_166__7), .B1 (nx66084)) ;
    dffr reg_ram_167__7 (.Q (ram_167__7), .QB (\$dummy [2022]), .D (nx51790), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51791 (.Y (nx51790), .A0 (ram_167__7), .A1 (nx65514), .S0 (
             nx63478)) ;
    dffr reg_ram_166__7 (.Q (ram_166__7), .QB (\$dummy [2023]), .D (nx51800), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51801 (.Y (nx51800), .A0 (ram_166__7), .A1 (nx65516), .S0 (
             nx63482)) ;
    nand04 ix20769 (.Y (nx20768), .A0 (nx63167), .A1 (nx63175), .A2 (nx63183), .A3 (
           nx63191)) ;
    aoi22 ix63168 (.Y (nx63167), .A0 (ram_168__7), .A1 (nx66088), .B0 (
          ram_169__7), .B1 (nx66092)) ;
    dffr reg_ram_168__7 (.Q (ram_168__7), .QB (\$dummy [2024]), .D (nx51780), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51781 (.Y (nx51780), .A0 (ram_168__7), .A1 (nx65516), .S0 (
             nx63474)) ;
    dffr reg_ram_169__7 (.Q (ram_169__7), .QB (\$dummy [2025]), .D (nx51770), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51771 (.Y (nx51770), .A0 (ram_169__7), .A1 (nx65516), .S0 (
             nx63470)) ;
    aoi22 ix63176 (.Y (nx63175), .A0 (ram_171__7), .A1 (nx66096), .B0 (
          ram_170__7), .B1 (nx66100)) ;
    dffr reg_ram_171__7 (.Q (ram_171__7), .QB (\$dummy [2026]), .D (nx51750), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51751 (.Y (nx51750), .A0 (ram_171__7), .A1 (nx65516), .S0 (
             nx63462)) ;
    dffr reg_ram_170__7 (.Q (ram_170__7), .QB (\$dummy [2027]), .D (nx51760), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51761 (.Y (nx51760), .A0 (ram_170__7), .A1 (nx65516), .S0 (
             nx63466)) ;
    aoi22 ix63184 (.Y (nx63183), .A0 (ram_172__7), .A1 (nx66104), .B0 (
          ram_173__7), .B1 (nx66108)) ;
    dffr reg_ram_172__7 (.Q (ram_172__7), .QB (\$dummy [2028]), .D (nx51740), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51741 (.Y (nx51740), .A0 (ram_172__7), .A1 (nx65516), .S0 (
             nx63458)) ;
    dffr reg_ram_173__7 (.Q (ram_173__7), .QB (\$dummy [2029]), .D (nx51730), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51731 (.Y (nx51730), .A0 (ram_173__7), .A1 (nx65516), .S0 (
             nx63454)) ;
    aoi22 ix63192 (.Y (nx63191), .A0 (ram_175__7), .A1 (nx66112), .B0 (
          ram_174__7), .B1 (nx66116)) ;
    dffr reg_ram_175__7 (.Q (ram_175__7), .QB (\$dummy [2030]), .D (nx51710), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51711 (.Y (nx51710), .A0 (ram_175__7), .A1 (nx65518), .S0 (
             nx63446)) ;
    dffr reg_ram_174__7 (.Q (ram_174__7), .QB (\$dummy [2031]), .D (nx51720), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51721 (.Y (nx51720), .A0 (ram_174__7), .A1 (nx65518), .S0 (
             nx63450)) ;
    oai21 ix63200 (.Y (nx63199), .A0 (nx20684), .A1 (nx20606), .B0 (nx66176)) ;
    nand04 ix20685 (.Y (nx20684), .A0 (nx63202), .A1 (nx63210), .A2 (nx63218), .A3 (
           nx63226)) ;
    aoi22 ix63203 (.Y (nx63202), .A0 (ram_176__7), .A1 (nx66056), .B0 (
          ram_177__7), .B1 (nx66060)) ;
    dffr reg_ram_176__7 (.Q (ram_176__7), .QB (\$dummy [2032]), .D (nx51700), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51701 (.Y (nx51700), .A0 (ram_176__7), .A1 (nx65518), .S0 (
             nx63436)) ;
    dffr reg_ram_177__7 (.Q (ram_177__7), .QB (\$dummy [2033]), .D (nx51690), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51691 (.Y (nx51690), .A0 (ram_177__7), .A1 (nx65518), .S0 (
             nx63426)) ;
    aoi22 ix63211 (.Y (nx63210), .A0 (ram_179__7), .A1 (nx66064), .B0 (
          ram_178__7), .B1 (nx66068)) ;
    dffr reg_ram_179__7 (.Q (ram_179__7), .QB (\$dummy [2034]), .D (nx51670), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51671 (.Y (nx51670), .A0 (ram_179__7), .A1 (nx65518), .S0 (
             nx63406)) ;
    dffr reg_ram_178__7 (.Q (ram_178__7), .QB (\$dummy [2035]), .D (nx51680), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51681 (.Y (nx51680), .A0 (ram_178__7), .A1 (nx65518), .S0 (
             nx63416)) ;
    aoi22 ix63219 (.Y (nx63218), .A0 (ram_180__7), .A1 (nx66072), .B0 (
          ram_181__7), .B1 (nx66076)) ;
    dffr reg_ram_180__7 (.Q (ram_180__7), .QB (\$dummy [2036]), .D (nx51660), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51661 (.Y (nx51660), .A0 (ram_180__7), .A1 (nx65518), .S0 (
             nx63396)) ;
    dffr reg_ram_181__7 (.Q (ram_181__7), .QB (\$dummy [2037]), .D (nx51650), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51651 (.Y (nx51650), .A0 (ram_181__7), .A1 (nx65520), .S0 (
             nx63386)) ;
    aoi22 ix63227 (.Y (nx63226), .A0 (ram_183__7), .A1 (nx66080), .B0 (
          ram_182__7), .B1 (nx66084)) ;
    dffr reg_ram_183__7 (.Q (ram_183__7), .QB (\$dummy [2038]), .D (nx51630), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51631 (.Y (nx51630), .A0 (ram_183__7), .A1 (nx65520), .S0 (
             nx63366)) ;
    dffr reg_ram_182__7 (.Q (ram_182__7), .QB (\$dummy [2039]), .D (nx51640), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51641 (.Y (nx51640), .A0 (ram_182__7), .A1 (nx65520), .S0 (
             nx63376)) ;
    nand04 ix20607 (.Y (nx20606), .A0 (nx63235), .A1 (nx63243), .A2 (nx63251), .A3 (
           nx63259)) ;
    aoi22 ix63236 (.Y (nx63235), .A0 (ram_184__7), .A1 (nx66088), .B0 (
          ram_185__7), .B1 (nx66092)) ;
    dffr reg_ram_184__7 (.Q (ram_184__7), .QB (\$dummy [2040]), .D (nx51620), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51621 (.Y (nx51620), .A0 (ram_184__7), .A1 (nx65520), .S0 (
             nx63356)) ;
    dffr reg_ram_185__7 (.Q (ram_185__7), .QB (\$dummy [2041]), .D (nx51610), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51611 (.Y (nx51610), .A0 (ram_185__7), .A1 (nx65520), .S0 (
             nx63346)) ;
    aoi22 ix63244 (.Y (nx63243), .A0 (ram_187__7), .A1 (nx66096), .B0 (
          ram_186__7), .B1 (nx66100)) ;
    dffr reg_ram_187__7 (.Q (ram_187__7), .QB (\$dummy [2042]), .D (nx51590), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51591 (.Y (nx51590), .A0 (ram_187__7), .A1 (nx65520), .S0 (
             nx63326)) ;
    dffr reg_ram_186__7 (.Q (ram_186__7), .QB (\$dummy [2043]), .D (nx51600), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51601 (.Y (nx51600), .A0 (ram_186__7), .A1 (nx65520), .S0 (
             nx63336)) ;
    aoi22 ix63252 (.Y (nx63251), .A0 (ram_188__7), .A1 (nx66104), .B0 (
          ram_189__7), .B1 (nx66108)) ;
    dffr reg_ram_188__7 (.Q (ram_188__7), .QB (\$dummy [2044]), .D (nx51580), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51581 (.Y (nx51580), .A0 (ram_188__7), .A1 (nx65522), .S0 (
             nx63316)) ;
    dffr reg_ram_189__7 (.Q (ram_189__7), .QB (\$dummy [2045]), .D (nx51570), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51571 (.Y (nx51570), .A0 (ram_189__7), .A1 (nx65522), .S0 (
             nx63306)) ;
    aoi22 ix63260 (.Y (nx63259), .A0 (ram_191__7), .A1 (nx66112), .B0 (
          ram_190__7), .B1 (nx66116)) ;
    dffr reg_ram_191__7 (.Q (ram_191__7), .QB (\$dummy [2046]), .D (nx51550), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51551 (.Y (nx51550), .A0 (ram_191__7), .A1 (nx65522), .S0 (
             nx63286)) ;
    dffr reg_ram_190__7 (.Q (ram_190__7), .QB (\$dummy [2047]), .D (nx51560), .CLK (
         clk), .R (rst)) ;
    mux21_ni ix51561 (.Y (nx51560), .A0 (ram_190__7), .A1 (nx65522), .S0 (
             nx63296)) ;
    buf02 ix63283 (.Y (nx63284), .A (nx32)) ;
    buf02 ix63285 (.Y (nx63286), .A (nx32)) ;
    buf02 ix63293 (.Y (nx63294), .A (nx54)) ;
    buf02 ix63295 (.Y (nx63296), .A (nx54)) ;
    buf02 ix63303 (.Y (nx63304), .A (nx78)) ;
    buf02 ix63305 (.Y (nx63306), .A (nx78)) ;
    buf02 ix63313 (.Y (nx63314), .A (nx98)) ;
    buf02 ix63315 (.Y (nx63316), .A (nx98)) ;
    buf02 ix63323 (.Y (nx63324), .A (nx124)) ;
    buf02 ix63325 (.Y (nx63326), .A (nx124)) ;
    buf02 ix63333 (.Y (nx63334), .A (nx142)) ;
    buf02 ix63335 (.Y (nx63336), .A (nx142)) ;
    buf02 ix63343 (.Y (nx63344), .A (nx162)) ;
    buf02 ix63345 (.Y (nx63346), .A (nx162)) ;
    buf02 ix63353 (.Y (nx63354), .A (nx180)) ;
    buf02 ix63355 (.Y (nx63356), .A (nx180)) ;
    buf02 ix63363 (.Y (nx63364), .A (nx208)) ;
    buf02 ix63365 (.Y (nx63366), .A (nx208)) ;
    buf02 ix63373 (.Y (nx63374), .A (nx226)) ;
    buf02 ix63375 (.Y (nx63376), .A (nx226)) ;
    buf02 ix63383 (.Y (nx63384), .A (nx246)) ;
    buf02 ix63385 (.Y (nx63386), .A (nx246)) ;
    buf02 ix63393 (.Y (nx63394), .A (nx264)) ;
    buf02 ix63395 (.Y (nx63396), .A (nx264)) ;
    buf02 ix63403 (.Y (nx63404), .A (nx288)) ;
    buf02 ix63405 (.Y (nx63406), .A (nx288)) ;
    buf02 ix63413 (.Y (nx63414), .A (nx306)) ;
    buf02 ix63415 (.Y (nx63416), .A (nx306)) ;
    buf02 ix63423 (.Y (nx63424), .A (nx326)) ;
    buf02 ix63425 (.Y (nx63426), .A (nx326)) ;
    buf02 ix63433 (.Y (nx63434), .A (nx344)) ;
    buf02 ix63435 (.Y (nx63436), .A (nx344)) ;
    buf02 ix63443 (.Y (nx63444), .A (nx378)) ;
    buf02 ix63445 (.Y (nx63446), .A (nx378)) ;
    buf02 ix63447 (.Y (nx63448), .A (nx394)) ;
    buf02 ix63449 (.Y (nx63450), .A (nx394)) ;
    buf02 ix63451 (.Y (nx63452), .A (nx412)) ;
    buf02 ix63453 (.Y (nx63454), .A (nx412)) ;
    buf02 ix63455 (.Y (nx63456), .A (nx428)) ;
    buf02 ix63457 (.Y (nx63458), .A (nx428)) ;
    buf02 ix63459 (.Y (nx63460), .A (nx448)) ;
    buf02 ix63461 (.Y (nx63462), .A (nx448)) ;
    buf02 ix63463 (.Y (nx63464), .A (nx464)) ;
    buf02 ix63465 (.Y (nx63466), .A (nx464)) ;
    buf02 ix63467 (.Y (nx63468), .A (nx482)) ;
    buf02 ix63469 (.Y (nx63470), .A (nx482)) ;
    buf02 ix63471 (.Y (nx63472), .A (nx498)) ;
    buf02 ix63473 (.Y (nx63474), .A (nx498)) ;
    buf02 ix63475 (.Y (nx63476), .A (nx520)) ;
    buf02 ix63477 (.Y (nx63478), .A (nx520)) ;
    buf02 ix63479 (.Y (nx63480), .A (nx536)) ;
    buf02 ix63481 (.Y (nx63482), .A (nx536)) ;
    buf02 ix63483 (.Y (nx63484), .A (nx554)) ;
    buf02 ix63485 (.Y (nx63486), .A (nx554)) ;
    buf02 ix63487 (.Y (nx63488), .A (nx570)) ;
    buf02 ix63489 (.Y (nx63490), .A (nx570)) ;
    buf02 ix63491 (.Y (nx63492), .A (nx590)) ;
    buf02 ix63493 (.Y (nx63494), .A (nx590)) ;
    buf02 ix63495 (.Y (nx63496), .A (nx606)) ;
    buf02 ix63497 (.Y (nx63498), .A (nx606)) ;
    buf02 ix63499 (.Y (nx63500), .A (nx624)) ;
    buf02 ix63501 (.Y (nx63502), .A (nx624)) ;
    buf02 ix63503 (.Y (nx63504), .A (nx640)) ;
    buf02 ix63505 (.Y (nx63506), .A (nx640)) ;
    buf02 ix63513 (.Y (nx63514), .A (nx676)) ;
    buf02 ix63515 (.Y (nx63516), .A (nx676)) ;
    buf02 ix63517 (.Y (nx63518), .A (nx692)) ;
    buf02 ix63519 (.Y (nx63520), .A (nx692)) ;
    buf02 ix63521 (.Y (nx63522), .A (nx710)) ;
    buf02 ix63523 (.Y (nx63524), .A (nx710)) ;
    buf02 ix63525 (.Y (nx63526), .A (nx726)) ;
    buf02 ix63527 (.Y (nx63528), .A (nx726)) ;
    buf02 ix63529 (.Y (nx63530), .A (nx746)) ;
    buf02 ix63531 (.Y (nx63532), .A (nx746)) ;
    buf02 ix63533 (.Y (nx63534), .A (nx762)) ;
    buf02 ix63535 (.Y (nx63536), .A (nx762)) ;
    buf02 ix63537 (.Y (nx63538), .A (nx780)) ;
    buf02 ix63539 (.Y (nx63540), .A (nx780)) ;
    buf02 ix63541 (.Y (nx63542), .A (nx796)) ;
    buf02 ix63543 (.Y (nx63544), .A (nx796)) ;
    buf02 ix63545 (.Y (nx63546), .A (nx818)) ;
    buf02 ix63547 (.Y (nx63548), .A (nx818)) ;
    buf02 ix63549 (.Y (nx63550), .A (nx834)) ;
    buf02 ix63551 (.Y (nx63552), .A (nx834)) ;
    buf02 ix63553 (.Y (nx63554), .A (nx852)) ;
    buf02 ix63555 (.Y (nx63556), .A (nx852)) ;
    buf02 ix63557 (.Y (nx63558), .A (nx868)) ;
    buf02 ix63559 (.Y (nx63560), .A (nx868)) ;
    buf02 ix63561 (.Y (nx63562), .A (nx888)) ;
    buf02 ix63563 (.Y (nx63564), .A (nx888)) ;
    buf02 ix63565 (.Y (nx63566), .A (nx904)) ;
    buf02 ix63567 (.Y (nx63568), .A (nx904)) ;
    buf02 ix63569 (.Y (nx63570), .A (nx922)) ;
    buf02 ix63571 (.Y (nx63572), .A (nx922)) ;
    buf02 ix63573 (.Y (nx63574), .A (nx938)) ;
    buf02 ix63575 (.Y (nx63576), .A (nx938)) ;
    buf02 ix63583 (.Y (nx63584), .A (nx970)) ;
    buf02 ix63585 (.Y (nx63586), .A (nx970)) ;
    buf02 ix63587 (.Y (nx63588), .A (nx986)) ;
    buf02 ix63589 (.Y (nx63590), .A (nx986)) ;
    buf02 ix63591 (.Y (nx63592), .A (nx1004)) ;
    buf02 ix63593 (.Y (nx63594), .A (nx1004)) ;
    buf02 ix63595 (.Y (nx63596), .A (nx1020)) ;
    buf02 ix63597 (.Y (nx63598), .A (nx1020)) ;
    buf02 ix63599 (.Y (nx63600), .A (nx1040)) ;
    buf02 ix63601 (.Y (nx63602), .A (nx1040)) ;
    buf02 ix63603 (.Y (nx63604), .A (nx1056)) ;
    buf02 ix63605 (.Y (nx63606), .A (nx1056)) ;
    buf02 ix63607 (.Y (nx63608), .A (nx1074)) ;
    buf02 ix63609 (.Y (nx63610), .A (nx1074)) ;
    buf02 ix63611 (.Y (nx63612), .A (nx1090)) ;
    buf02 ix63613 (.Y (nx63614), .A (nx1090)) ;
    buf02 ix63615 (.Y (nx63616), .A (nx1112)) ;
    buf02 ix63617 (.Y (nx63618), .A (nx1112)) ;
    buf02 ix63619 (.Y (nx63620), .A (nx1128)) ;
    buf02 ix63621 (.Y (nx63622), .A (nx1128)) ;
    buf02 ix63623 (.Y (nx63624), .A (nx1146)) ;
    buf02 ix63625 (.Y (nx63626), .A (nx1146)) ;
    buf02 ix63627 (.Y (nx63628), .A (nx1162)) ;
    buf02 ix63629 (.Y (nx63630), .A (nx1162)) ;
    buf02 ix63631 (.Y (nx63632), .A (nx1182)) ;
    buf02 ix63633 (.Y (nx63634), .A (nx1182)) ;
    buf02 ix63635 (.Y (nx63636), .A (nx1198)) ;
    buf02 ix63637 (.Y (nx63638), .A (nx1198)) ;
    buf02 ix63639 (.Y (nx63640), .A (nx1216)) ;
    buf02 ix63641 (.Y (nx63642), .A (nx1216)) ;
    buf02 ix63643 (.Y (nx63644), .A (nx1232)) ;
    buf02 ix63645 (.Y (nx63646), .A (nx1232)) ;
    buf02 ix63653 (.Y (nx63654), .A (nx1270)) ;
    buf02 ix63655 (.Y (nx63656), .A (nx1270)) ;
    buf02 ix63657 (.Y (nx63658), .A (nx1286)) ;
    buf02 ix63659 (.Y (nx63660), .A (nx1286)) ;
    buf02 ix63661 (.Y (nx63662), .A (nx1304)) ;
    buf02 ix63663 (.Y (nx63664), .A (nx1304)) ;
    buf02 ix63665 (.Y (nx63666), .A (nx1320)) ;
    buf02 ix63667 (.Y (nx63668), .A (nx1320)) ;
    buf02 ix63669 (.Y (nx63670), .A (nx1340)) ;
    buf02 ix63671 (.Y (nx63672), .A (nx1340)) ;
    buf02 ix63673 (.Y (nx63674), .A (nx1356)) ;
    buf02 ix63675 (.Y (nx63676), .A (nx1356)) ;
    buf02 ix63677 (.Y (nx63678), .A (nx1374)) ;
    buf02 ix63679 (.Y (nx63680), .A (nx1374)) ;
    buf02 ix63681 (.Y (nx63682), .A (nx1390)) ;
    buf02 ix63683 (.Y (nx63684), .A (nx1390)) ;
    buf02 ix63685 (.Y (nx63686), .A (nx1412)) ;
    buf02 ix63687 (.Y (nx63688), .A (nx1412)) ;
    buf02 ix63689 (.Y (nx63690), .A (nx1428)) ;
    buf02 ix63691 (.Y (nx63692), .A (nx1428)) ;
    buf02 ix63693 (.Y (nx63694), .A (nx1446)) ;
    buf02 ix63695 (.Y (nx63696), .A (nx1446)) ;
    buf02 ix63697 (.Y (nx63698), .A (nx1462)) ;
    buf02 ix63699 (.Y (nx63700), .A (nx1462)) ;
    buf02 ix63701 (.Y (nx63702), .A (nx1482)) ;
    buf02 ix63703 (.Y (nx63704), .A (nx1482)) ;
    buf02 ix63705 (.Y (nx63706), .A (nx1498)) ;
    buf02 ix63707 (.Y (nx63708), .A (nx1498)) ;
    buf02 ix63709 (.Y (nx63710), .A (nx1516)) ;
    buf02 ix63711 (.Y (nx63712), .A (nx1516)) ;
    buf02 ix63713 (.Y (nx63714), .A (nx1532)) ;
    buf02 ix63715 (.Y (nx63716), .A (nx1532)) ;
    buf02 ix63723 (.Y (nx63724), .A (nx1562)) ;
    buf02 ix63725 (.Y (nx63726), .A (nx1562)) ;
    buf02 ix63727 (.Y (nx63728), .A (nx1578)) ;
    buf02 ix63729 (.Y (nx63730), .A (nx1578)) ;
    buf02 ix63731 (.Y (nx63732), .A (nx1596)) ;
    buf02 ix63733 (.Y (nx63734), .A (nx1596)) ;
    buf02 ix63735 (.Y (nx63736), .A (nx1612)) ;
    buf02 ix63737 (.Y (nx63738), .A (nx1612)) ;
    buf02 ix63739 (.Y (nx63740), .A (nx1632)) ;
    buf02 ix63741 (.Y (nx63742), .A (nx1632)) ;
    buf02 ix63743 (.Y (nx63744), .A (nx1648)) ;
    buf02 ix63745 (.Y (nx63746), .A (nx1648)) ;
    buf02 ix63747 (.Y (nx63748), .A (nx1666)) ;
    buf02 ix63749 (.Y (nx63750), .A (nx1666)) ;
    buf02 ix63751 (.Y (nx63752), .A (nx1682)) ;
    buf02 ix63753 (.Y (nx63754), .A (nx1682)) ;
    buf02 ix63755 (.Y (nx63756), .A (nx1704)) ;
    buf02 ix63757 (.Y (nx63758), .A (nx1704)) ;
    buf02 ix63759 (.Y (nx63760), .A (nx1720)) ;
    buf02 ix63761 (.Y (nx63762), .A (nx1720)) ;
    buf02 ix63763 (.Y (nx63764), .A (nx1738)) ;
    buf02 ix63765 (.Y (nx63766), .A (nx1738)) ;
    buf02 ix63767 (.Y (nx63768), .A (nx1754)) ;
    buf02 ix63769 (.Y (nx63770), .A (nx1754)) ;
    buf02 ix63771 (.Y (nx63772), .A (nx1774)) ;
    buf02 ix63773 (.Y (nx63774), .A (nx1774)) ;
    buf02 ix63775 (.Y (nx63776), .A (nx1790)) ;
    buf02 ix63777 (.Y (nx63778), .A (nx1790)) ;
    buf02 ix63779 (.Y (nx63780), .A (nx1808)) ;
    buf02 ix63781 (.Y (nx63782), .A (nx1808)) ;
    buf02 ix63783 (.Y (nx63784), .A (nx1824)) ;
    buf02 ix63785 (.Y (nx63786), .A (nx1824)) ;
    buf02 ix63793 (.Y (nx63794), .A (nx2150)) ;
    buf02 ix63795 (.Y (nx63796), .A (nx2150)) ;
    buf02 ix63797 (.Y (nx63798), .A (nx2166)) ;
    buf02 ix63799 (.Y (nx63800), .A (nx2166)) ;
    buf02 ix63801 (.Y (nx63802), .A (nx2184)) ;
    buf02 ix63803 (.Y (nx63804), .A (nx2184)) ;
    buf02 ix63805 (.Y (nx63806), .A (nx2200)) ;
    buf02 ix63807 (.Y (nx63808), .A (nx2200)) ;
    buf02 ix63809 (.Y (nx63810), .A (nx2220)) ;
    buf02 ix63811 (.Y (nx63812), .A (nx2220)) ;
    buf02 ix63813 (.Y (nx63814), .A (nx2236)) ;
    buf02 ix63815 (.Y (nx63816), .A (nx2236)) ;
    buf02 ix63817 (.Y (nx63818), .A (nx2254)) ;
    buf02 ix63819 (.Y (nx63820), .A (nx2254)) ;
    buf02 ix63821 (.Y (nx63822), .A (nx2270)) ;
    buf02 ix63823 (.Y (nx63824), .A (nx2270)) ;
    buf02 ix63825 (.Y (nx63826), .A (nx2292)) ;
    buf02 ix63827 (.Y (nx63828), .A (nx2292)) ;
    buf02 ix63829 (.Y (nx63830), .A (nx2308)) ;
    buf02 ix63831 (.Y (nx63832), .A (nx2308)) ;
    buf02 ix63833 (.Y (nx63834), .A (nx2326)) ;
    buf02 ix63835 (.Y (nx63836), .A (nx2326)) ;
    buf02 ix63837 (.Y (nx63838), .A (nx2342)) ;
    buf02 ix63839 (.Y (nx63840), .A (nx2342)) ;
    buf02 ix63841 (.Y (nx63842), .A (nx2362)) ;
    buf02 ix63843 (.Y (nx63844), .A (nx2362)) ;
    buf02 ix63845 (.Y (nx63846), .A (nx2378)) ;
    buf02 ix63847 (.Y (nx63848), .A (nx2378)) ;
    buf02 ix63849 (.Y (nx63850), .A (nx2396)) ;
    buf02 ix63851 (.Y (nx63852), .A (nx2396)) ;
    buf02 ix63853 (.Y (nx63854), .A (nx2412)) ;
    buf02 ix63855 (.Y (nx63856), .A (nx2412)) ;
    buf02 ix63863 (.Y (nx63864), .A (nx2448)) ;
    buf02 ix63865 (.Y (nx63866), .A (nx2448)) ;
    buf02 ix63867 (.Y (nx63868), .A (nx2464)) ;
    buf02 ix63869 (.Y (nx63870), .A (nx2464)) ;
    buf02 ix63871 (.Y (nx63872), .A (nx2482)) ;
    buf02 ix63873 (.Y (nx63874), .A (nx2482)) ;
    buf02 ix63875 (.Y (nx63876), .A (nx2498)) ;
    buf02 ix63877 (.Y (nx63878), .A (nx2498)) ;
    buf02 ix63879 (.Y (nx63880), .A (nx2518)) ;
    buf02 ix63881 (.Y (nx63882), .A (nx2518)) ;
    buf02 ix63883 (.Y (nx63884), .A (nx2534)) ;
    buf02 ix63885 (.Y (nx63886), .A (nx2534)) ;
    buf02 ix63887 (.Y (nx63888), .A (nx2552)) ;
    buf02 ix63889 (.Y (nx63890), .A (nx2552)) ;
    buf02 ix63891 (.Y (nx63892), .A (nx2568)) ;
    buf02 ix63893 (.Y (nx63894), .A (nx2568)) ;
    buf02 ix63895 (.Y (nx63896), .A (nx2590)) ;
    buf02 ix63897 (.Y (nx63898), .A (nx2590)) ;
    buf02 ix63899 (.Y (nx63900), .A (nx2606)) ;
    buf02 ix63901 (.Y (nx63902), .A (nx2606)) ;
    buf02 ix63903 (.Y (nx63904), .A (nx2624)) ;
    buf02 ix63905 (.Y (nx63906), .A (nx2624)) ;
    buf02 ix63907 (.Y (nx63908), .A (nx2640)) ;
    buf02 ix63909 (.Y (nx63910), .A (nx2640)) ;
    buf02 ix63911 (.Y (nx63912), .A (nx2660)) ;
    buf02 ix63913 (.Y (nx63914), .A (nx2660)) ;
    buf02 ix63915 (.Y (nx63916), .A (nx2676)) ;
    buf02 ix63917 (.Y (nx63918), .A (nx2676)) ;
    buf02 ix63919 (.Y (nx63920), .A (nx2694)) ;
    buf02 ix63921 (.Y (nx63922), .A (nx2694)) ;
    buf02 ix63923 (.Y (nx63924), .A (nx2710)) ;
    buf02 ix63925 (.Y (nx63926), .A (nx2710)) ;
    buf02 ix63933 (.Y (nx63934), .A (nx2740)) ;
    buf02 ix63935 (.Y (nx63936), .A (nx2740)) ;
    buf02 ix63937 (.Y (nx63938), .A (nx2756)) ;
    buf02 ix63939 (.Y (nx63940), .A (nx2756)) ;
    buf02 ix63941 (.Y (nx63942), .A (nx2774)) ;
    buf02 ix63943 (.Y (nx63944), .A (nx2774)) ;
    buf02 ix63945 (.Y (nx63946), .A (nx2790)) ;
    buf02 ix63947 (.Y (nx63948), .A (nx2790)) ;
    buf02 ix63949 (.Y (nx63950), .A (nx2810)) ;
    buf02 ix63951 (.Y (nx63952), .A (nx2810)) ;
    buf02 ix63953 (.Y (nx63954), .A (nx2826)) ;
    buf02 ix63955 (.Y (nx63956), .A (nx2826)) ;
    buf02 ix63957 (.Y (nx63958), .A (nx2844)) ;
    buf02 ix63959 (.Y (nx63960), .A (nx2844)) ;
    buf02 ix63961 (.Y (nx63962), .A (nx2860)) ;
    buf02 ix63963 (.Y (nx63964), .A (nx2860)) ;
    buf02 ix63965 (.Y (nx63966), .A (nx2882)) ;
    buf02 ix63967 (.Y (nx63968), .A (nx2882)) ;
    buf02 ix63969 (.Y (nx63970), .A (nx2898)) ;
    buf02 ix63971 (.Y (nx63972), .A (nx2898)) ;
    buf02 ix63973 (.Y (nx63974), .A (nx2916)) ;
    buf02 ix63975 (.Y (nx63976), .A (nx2916)) ;
    buf02 ix63977 (.Y (nx63978), .A (nx2932)) ;
    buf02 ix63979 (.Y (nx63980), .A (nx2932)) ;
    buf02 ix63981 (.Y (nx63982), .A (nx2952)) ;
    buf02 ix63983 (.Y (nx63984), .A (nx2952)) ;
    buf02 ix63985 (.Y (nx63986), .A (nx2968)) ;
    buf02 ix63987 (.Y (nx63988), .A (nx2968)) ;
    buf02 ix63989 (.Y (nx63990), .A (nx2986)) ;
    buf02 ix63991 (.Y (nx63992), .A (nx2986)) ;
    buf02 ix63993 (.Y (nx63994), .A (nx3002)) ;
    buf02 ix63995 (.Y (nx63996), .A (nx3002)) ;
    buf02 ix64003 (.Y (nx64004), .A (nx3034)) ;
    buf02 ix64005 (.Y (nx64006), .A (nx3034)) ;
    buf02 ix64007 (.Y (nx64008), .A (nx3050)) ;
    buf02 ix64009 (.Y (nx64010), .A (nx3050)) ;
    buf02 ix64011 (.Y (nx64012), .A (nx3068)) ;
    buf02 ix64013 (.Y (nx64014), .A (nx3068)) ;
    buf02 ix64015 (.Y (nx64016), .A (nx3084)) ;
    buf02 ix64017 (.Y (nx64018), .A (nx3084)) ;
    buf02 ix64019 (.Y (nx64020), .A (nx3104)) ;
    buf02 ix64021 (.Y (nx64022), .A (nx3104)) ;
    buf02 ix64023 (.Y (nx64024), .A (nx3120)) ;
    buf02 ix64025 (.Y (nx64026), .A (nx3120)) ;
    buf02 ix64027 (.Y (nx64028), .A (nx3138)) ;
    buf02 ix64029 (.Y (nx64030), .A (nx3138)) ;
    buf02 ix64031 (.Y (nx64032), .A (nx3154)) ;
    buf02 ix64033 (.Y (nx64034), .A (nx3154)) ;
    buf02 ix64035 (.Y (nx64036), .A (nx3176)) ;
    buf02 ix64037 (.Y (nx64038), .A (nx3176)) ;
    buf02 ix64039 (.Y (nx64040), .A (nx3192)) ;
    buf02 ix64041 (.Y (nx64042), .A (nx3192)) ;
    buf02 ix64043 (.Y (nx64044), .A (nx3210)) ;
    buf02 ix64045 (.Y (nx64046), .A (nx3210)) ;
    buf02 ix64047 (.Y (nx64048), .A (nx3226)) ;
    buf02 ix64049 (.Y (nx64050), .A (nx3226)) ;
    buf02 ix64051 (.Y (nx64052), .A (nx3246)) ;
    buf02 ix64053 (.Y (nx64054), .A (nx3246)) ;
    buf02 ix64055 (.Y (nx64056), .A (nx3262)) ;
    buf02 ix64057 (.Y (nx64058), .A (nx3262)) ;
    buf02 ix64059 (.Y (nx64060), .A (nx3280)) ;
    buf02 ix64061 (.Y (nx64062), .A (nx3280)) ;
    buf02 ix64063 (.Y (nx64064), .A (nx3296)) ;
    buf02 ix64065 (.Y (nx64066), .A (nx3296)) ;
    buf02 ix64073 (.Y (nx64074), .A (nx3326)) ;
    buf02 ix64075 (.Y (nx64076), .A (nx3326)) ;
    buf02 ix64077 (.Y (nx64078), .A (nx3342)) ;
    buf02 ix64079 (.Y (nx64080), .A (nx3342)) ;
    buf02 ix64081 (.Y (nx64082), .A (nx3360)) ;
    buf02 ix64083 (.Y (nx64084), .A (nx3360)) ;
    buf02 ix64085 (.Y (nx64086), .A (nx3376)) ;
    buf02 ix64087 (.Y (nx64088), .A (nx3376)) ;
    buf02 ix64089 (.Y (nx64090), .A (nx3396)) ;
    buf02 ix64091 (.Y (nx64092), .A (nx3396)) ;
    buf02 ix64093 (.Y (nx64094), .A (nx3412)) ;
    buf02 ix64095 (.Y (nx64096), .A (nx3412)) ;
    buf02 ix64097 (.Y (nx64098), .A (nx3430)) ;
    buf02 ix64099 (.Y (nx64100), .A (nx3430)) ;
    buf02 ix64101 (.Y (nx64102), .A (nx3446)) ;
    buf02 ix64103 (.Y (nx64104), .A (nx3446)) ;
    buf02 ix64105 (.Y (nx64106), .A (nx3468)) ;
    buf02 ix64107 (.Y (nx64108), .A (nx3468)) ;
    buf02 ix64109 (.Y (nx64110), .A (nx3484)) ;
    buf02 ix64111 (.Y (nx64112), .A (nx3484)) ;
    buf02 ix64113 (.Y (nx64114), .A (nx3502)) ;
    buf02 ix64115 (.Y (nx64116), .A (nx3502)) ;
    buf02 ix64117 (.Y (nx64118), .A (nx3518)) ;
    buf02 ix64119 (.Y (nx64120), .A (nx3518)) ;
    buf02 ix64121 (.Y (nx64122), .A (nx3538)) ;
    buf02 ix64123 (.Y (nx64124), .A (nx3538)) ;
    buf02 ix64125 (.Y (nx64126), .A (nx3554)) ;
    buf02 ix64127 (.Y (nx64128), .A (nx3554)) ;
    buf02 ix64129 (.Y (nx64130), .A (nx3572)) ;
    buf02 ix64131 (.Y (nx64132), .A (nx3572)) ;
    buf02 ix64133 (.Y (nx64134), .A (nx3588)) ;
    buf02 ix64135 (.Y (nx64136), .A (nx3588)) ;
    buf02 ix64143 (.Y (nx64144), .A (nx3628)) ;
    buf02 ix64145 (.Y (nx64146), .A (nx3628)) ;
    buf02 ix64147 (.Y (nx64148), .A (nx3644)) ;
    buf02 ix64149 (.Y (nx64150), .A (nx3644)) ;
    buf02 ix64151 (.Y (nx64152), .A (nx3662)) ;
    buf02 ix64153 (.Y (nx64154), .A (nx3662)) ;
    buf02 ix64155 (.Y (nx64156), .A (nx3678)) ;
    buf02 ix64157 (.Y (nx64158), .A (nx3678)) ;
    buf02 ix64159 (.Y (nx64160), .A (nx3698)) ;
    buf02 ix64161 (.Y (nx64162), .A (nx3698)) ;
    buf02 ix64163 (.Y (nx64164), .A (nx3714)) ;
    buf02 ix64165 (.Y (nx64166), .A (nx3714)) ;
    buf02 ix64167 (.Y (nx64168), .A (nx3732)) ;
    buf02 ix64169 (.Y (nx64170), .A (nx3732)) ;
    buf02 ix64171 (.Y (nx64172), .A (nx3748)) ;
    buf02 ix64173 (.Y (nx64174), .A (nx3748)) ;
    buf02 ix64175 (.Y (nx64176), .A (nx3770)) ;
    buf02 ix64177 (.Y (nx64178), .A (nx3770)) ;
    buf02 ix64179 (.Y (nx64180), .A (nx3786)) ;
    buf02 ix64181 (.Y (nx64182), .A (nx3786)) ;
    buf02 ix64183 (.Y (nx64184), .A (nx3804)) ;
    buf02 ix64185 (.Y (nx64186), .A (nx3804)) ;
    buf02 ix64187 (.Y (nx64188), .A (nx3820)) ;
    buf02 ix64189 (.Y (nx64190), .A (nx3820)) ;
    buf02 ix64191 (.Y (nx64192), .A (nx3840)) ;
    buf02 ix64193 (.Y (nx64194), .A (nx3840)) ;
    buf02 ix64195 (.Y (nx64196), .A (nx3856)) ;
    buf02 ix64197 (.Y (nx64198), .A (nx3856)) ;
    buf02 ix64199 (.Y (nx64200), .A (nx3874)) ;
    buf02 ix64201 (.Y (nx64202), .A (nx3874)) ;
    buf02 ix64203 (.Y (nx64204), .A (nx3890)) ;
    buf02 ix64205 (.Y (nx64206), .A (nx3890)) ;
    buf02 ix64213 (.Y (nx64214), .A (nx3920)) ;
    buf02 ix64215 (.Y (nx64216), .A (nx3920)) ;
    buf02 ix64217 (.Y (nx64218), .A (nx3936)) ;
    buf02 ix64219 (.Y (nx64220), .A (nx3936)) ;
    buf02 ix64221 (.Y (nx64222), .A (nx3954)) ;
    buf02 ix64223 (.Y (nx64224), .A (nx3954)) ;
    buf02 ix64225 (.Y (nx64226), .A (nx3970)) ;
    buf02 ix64227 (.Y (nx64228), .A (nx3970)) ;
    buf02 ix64229 (.Y (nx64230), .A (nx3990)) ;
    buf02 ix64231 (.Y (nx64232), .A (nx3990)) ;
    buf02 ix64233 (.Y (nx64234), .A (nx4006)) ;
    buf02 ix64235 (.Y (nx64236), .A (nx4006)) ;
    buf02 ix64237 (.Y (nx64238), .A (nx4024)) ;
    buf02 ix64239 (.Y (nx64240), .A (nx4024)) ;
    buf02 ix64241 (.Y (nx64242), .A (nx4040)) ;
    buf02 ix64243 (.Y (nx64244), .A (nx4040)) ;
    buf02 ix64245 (.Y (nx64246), .A (nx4062)) ;
    buf02 ix64247 (.Y (nx64248), .A (nx4062)) ;
    buf02 ix64249 (.Y (nx64250), .A (nx4078)) ;
    buf02 ix64251 (.Y (nx64252), .A (nx4078)) ;
    buf02 ix64253 (.Y (nx64254), .A (nx4096)) ;
    buf02 ix64255 (.Y (nx64256), .A (nx4096)) ;
    buf02 ix64257 (.Y (nx64258), .A (nx4112)) ;
    buf02 ix64259 (.Y (nx64260), .A (nx4112)) ;
    buf02 ix64261 (.Y (nx64262), .A (nx4132)) ;
    buf02 ix64263 (.Y (nx64264), .A (nx4132)) ;
    buf02 ix64265 (.Y (nx64266), .A (nx4148)) ;
    buf02 ix64267 (.Y (nx64268), .A (nx4148)) ;
    buf02 ix64269 (.Y (nx64270), .A (nx4166)) ;
    buf02 ix64271 (.Y (nx64272), .A (nx4166)) ;
    buf02 ix64273 (.Y (nx64274), .A (nx4182)) ;
    buf02 ix64275 (.Y (nx64276), .A (nx4182)) ;
    buf02 ix64283 (.Y (nx64284), .A (nx4214)) ;
    buf02 ix64285 (.Y (nx64286), .A (nx4214)) ;
    buf02 ix64287 (.Y (nx64288), .A (nx4230)) ;
    buf02 ix64289 (.Y (nx64290), .A (nx4230)) ;
    buf02 ix64291 (.Y (nx64292), .A (nx4248)) ;
    buf02 ix64293 (.Y (nx64294), .A (nx4248)) ;
    buf02 ix64295 (.Y (nx64296), .A (nx4264)) ;
    buf02 ix64297 (.Y (nx64298), .A (nx4264)) ;
    buf02 ix64299 (.Y (nx64300), .A (nx4284)) ;
    buf02 ix64301 (.Y (nx64302), .A (nx4284)) ;
    buf02 ix64303 (.Y (nx64304), .A (nx4300)) ;
    buf02 ix64305 (.Y (nx64306), .A (nx4300)) ;
    buf02 ix64307 (.Y (nx64308), .A (nx4318)) ;
    buf02 ix64309 (.Y (nx64310), .A (nx4318)) ;
    buf02 ix64311 (.Y (nx64312), .A (nx4334)) ;
    buf02 ix64313 (.Y (nx64314), .A (nx4334)) ;
    buf02 ix64315 (.Y (nx64316), .A (nx4356)) ;
    buf02 ix64317 (.Y (nx64318), .A (nx4356)) ;
    buf02 ix64319 (.Y (nx64320), .A (nx4372)) ;
    buf02 ix64321 (.Y (nx64322), .A (nx4372)) ;
    buf02 ix64323 (.Y (nx64324), .A (nx4390)) ;
    buf02 ix64325 (.Y (nx64326), .A (nx4390)) ;
    buf02 ix64327 (.Y (nx64328), .A (nx4406)) ;
    buf02 ix64329 (.Y (nx64330), .A (nx4406)) ;
    buf02 ix64331 (.Y (nx64332), .A (nx4426)) ;
    buf02 ix64333 (.Y (nx64334), .A (nx4426)) ;
    buf02 ix64335 (.Y (nx64336), .A (nx4442)) ;
    buf02 ix64337 (.Y (nx64338), .A (nx4442)) ;
    buf02 ix64339 (.Y (nx64340), .A (nx4460)) ;
    buf02 ix64341 (.Y (nx64342), .A (nx4460)) ;
    buf02 ix64343 (.Y (nx64344), .A (nx4476)) ;
    buf02 ix64345 (.Y (nx64346), .A (nx4476)) ;
    buf02 ix64353 (.Y (nx64354), .A (nx4506)) ;
    buf02 ix64355 (.Y (nx64356), .A (nx4506)) ;
    buf02 ix64357 (.Y (nx64358), .A (nx4522)) ;
    buf02 ix64359 (.Y (nx64360), .A (nx4522)) ;
    buf02 ix64361 (.Y (nx64362), .A (nx4540)) ;
    buf02 ix64363 (.Y (nx64364), .A (nx4540)) ;
    buf02 ix64365 (.Y (nx64366), .A (nx4556)) ;
    buf02 ix64367 (.Y (nx64368), .A (nx4556)) ;
    buf02 ix64369 (.Y (nx64370), .A (nx4576)) ;
    buf02 ix64371 (.Y (nx64372), .A (nx4576)) ;
    buf02 ix64373 (.Y (nx64374), .A (nx4592)) ;
    buf02 ix64375 (.Y (nx64376), .A (nx4592)) ;
    buf02 ix64377 (.Y (nx64378), .A (nx4610)) ;
    buf02 ix64379 (.Y (nx64380), .A (nx4610)) ;
    buf02 ix64381 (.Y (nx64382), .A (nx4626)) ;
    buf02 ix64383 (.Y (nx64384), .A (nx4626)) ;
    buf02 ix64385 (.Y (nx64386), .A (nx4648)) ;
    buf02 ix64387 (.Y (nx64388), .A (nx4648)) ;
    buf02 ix64389 (.Y (nx64390), .A (nx4664)) ;
    buf02 ix64391 (.Y (nx64392), .A (nx4664)) ;
    buf02 ix64393 (.Y (nx64394), .A (nx4682)) ;
    buf02 ix64395 (.Y (nx64396), .A (nx4682)) ;
    buf02 ix64397 (.Y (nx64398), .A (nx4698)) ;
    buf02 ix64399 (.Y (nx64400), .A (nx4698)) ;
    buf02 ix64401 (.Y (nx64402), .A (nx4718)) ;
    buf02 ix64403 (.Y (nx64404), .A (nx4718)) ;
    buf02 ix64405 (.Y (nx64406), .A (nx4734)) ;
    buf02 ix64407 (.Y (nx64408), .A (nx4734)) ;
    buf02 ix64409 (.Y (nx64410), .A (nx4752)) ;
    buf02 ix64411 (.Y (nx64412), .A (nx4752)) ;
    buf02 ix64413 (.Y (nx64414), .A (nx4768)) ;
    buf02 ix64415 (.Y (nx64416), .A (nx4768)) ;
    inv02 ix64487 (.Y (nx64488), .A (nx65324)) ;
    inv02 ix64489 (.Y (nx64490), .A (nx65324)) ;
    inv02 ix64491 (.Y (nx64492), .A (nx65324)) ;
    inv02 ix64493 (.Y (nx64494), .A (nx65324)) ;
    inv02 ix64495 (.Y (nx64496), .A (nx65324)) ;
    inv02 ix64497 (.Y (nx64498), .A (nx65324)) ;
    inv02 ix64499 (.Y (nx64500), .A (nx65324)) ;
    inv02 ix64501 (.Y (nx64502), .A (nx65326)) ;
    inv02 ix64503 (.Y (nx64504), .A (nx65326)) ;
    inv02 ix64505 (.Y (nx64506), .A (nx65326)) ;
    inv02 ix64507 (.Y (nx64508), .A (nx65326)) ;
    inv02 ix64509 (.Y (nx64510), .A (nx65326)) ;
    inv02 ix64511 (.Y (nx64512), .A (nx65326)) ;
    inv02 ix64513 (.Y (nx64514), .A (nx65326)) ;
    inv02 ix64515 (.Y (nx64516), .A (nx65328)) ;
    inv02 ix64517 (.Y (nx64518), .A (nx65328)) ;
    inv02 ix64519 (.Y (nx64520), .A (nx65328)) ;
    inv02 ix64521 (.Y (nx64522), .A (nx65328)) ;
    inv02 ix64523 (.Y (nx64524), .A (nx65328)) ;
    inv02 ix64525 (.Y (nx64526), .A (nx318)) ;
    inv02 ix64527 (.Y (nx64528), .A (nx65318)) ;
    inv02 ix64529 (.Y (nx64530), .A (nx65318)) ;
    inv02 ix64531 (.Y (nx64532), .A (nx65318)) ;
    inv02 ix64533 (.Y (nx64534), .A (nx65318)) ;
    inv02 ix64535 (.Y (nx64536), .A (nx65318)) ;
    inv02 ix64537 (.Y (nx64538), .A (nx65318)) ;
    inv02 ix64539 (.Y (nx64540), .A (nx65318)) ;
    inv02 ix64541 (.Y (nx64542), .A (nx65320)) ;
    inv02 ix64543 (.Y (nx64544), .A (nx65320)) ;
    inv02 ix64545 (.Y (nx64546), .A (nx65320)) ;
    inv02 ix64547 (.Y (nx64548), .A (nx65320)) ;
    inv02 ix64549 (.Y (nx64550), .A (nx65320)) ;
    inv02 ix64551 (.Y (nx64552), .A (nx65320)) ;
    inv02 ix64553 (.Y (nx64554), .A (nx65320)) ;
    inv02 ix64555 (.Y (nx64556), .A (nx65322)) ;
    inv02 ix64557 (.Y (nx64558), .A (nx65322)) ;
    inv02 ix64559 (.Y (nx64560), .A (nx65322)) ;
    inv02 ix64561 (.Y (nx64562), .A (nx65322)) ;
    inv02 ix64563 (.Y (nx64564), .A (nx280)) ;
    inv02 ix64565 (.Y (nx64566), .A (nx65306)) ;
    inv02 ix64567 (.Y (nx64568), .A (nx65306)) ;
    inv02 ix64569 (.Y (nx64570), .A (nx65306)) ;
    inv02 ix64571 (.Y (nx64572), .A (nx65306)) ;
    inv02 ix64573 (.Y (nx64574), .A (nx65306)) ;
    inv02 ix64575 (.Y (nx64576), .A (nx65306)) ;
    inv02 ix64577 (.Y (nx64578), .A (nx65306)) ;
    inv02 ix64579 (.Y (nx64580), .A (nx65308)) ;
    inv02 ix64581 (.Y (nx64582), .A (nx65308)) ;
    inv02 ix64583 (.Y (nx64584), .A (nx65308)) ;
    inv02 ix64585 (.Y (nx64586), .A (nx65308)) ;
    inv02 ix64587 (.Y (nx64588), .A (nx65308)) ;
    inv02 ix64589 (.Y (nx64590), .A (nx65308)) ;
    inv02 ix64591 (.Y (nx64592), .A (nx65308)) ;
    inv02 ix64593 (.Y (nx64594), .A (nx65310)) ;
    inv02 ix64595 (.Y (nx64596), .A (nx65310)) ;
    inv02 ix64597 (.Y (nx64598), .A (nx65310)) ;
    inv02 ix64599 (.Y (nx64600), .A (nx65310)) ;
    inv02 ix64601 (.Y (nx64602), .A (nx298)) ;
    inv02 ix64603 (.Y (nx64604), .A (nx65312)) ;
    inv02 ix64605 (.Y (nx64606), .A (nx65312)) ;
    inv02 ix64607 (.Y (nx64608), .A (nx65312)) ;
    inv02 ix64609 (.Y (nx64610), .A (nx65312)) ;
    inv02 ix64611 (.Y (nx64612), .A (nx65312)) ;
    inv02 ix64613 (.Y (nx64614), .A (nx65312)) ;
    inv02 ix64615 (.Y (nx64616), .A (nx65312)) ;
    inv02 ix64617 (.Y (nx64618), .A (nx65314)) ;
    inv02 ix64619 (.Y (nx64620), .A (nx65314)) ;
    inv02 ix64621 (.Y (nx64622), .A (nx65314)) ;
    inv02 ix64623 (.Y (nx64624), .A (nx65314)) ;
    inv02 ix64625 (.Y (nx64626), .A (nx65314)) ;
    inv02 ix64627 (.Y (nx64628), .A (nx65314)) ;
    inv02 ix64629 (.Y (nx64630), .A (nx65314)) ;
    inv02 ix64631 (.Y (nx64632), .A (nx65316)) ;
    inv02 ix64633 (.Y (nx64634), .A (nx65316)) ;
    inv02 ix64635 (.Y (nx64636), .A (nx65316)) ;
    inv02 ix64637 (.Y (nx64638), .A (nx65316)) ;
    inv02 ix64639 (.Y (nx64640), .A (nx256)) ;
    inv02 ix64641 (.Y (nx64642), .A (nx65300)) ;
    inv02 ix64643 (.Y (nx64644), .A (nx65300)) ;
    inv02 ix64645 (.Y (nx64646), .A (nx65300)) ;
    inv02 ix64647 (.Y (nx64648), .A (nx65300)) ;
    inv02 ix64649 (.Y (nx64650), .A (nx65300)) ;
    inv02 ix64651 (.Y (nx64652), .A (nx65300)) ;
    inv02 ix64653 (.Y (nx64654), .A (nx65300)) ;
    inv02 ix64655 (.Y (nx64656), .A (nx65302)) ;
    inv02 ix64657 (.Y (nx64658), .A (nx65302)) ;
    inv02 ix64659 (.Y (nx64660), .A (nx65302)) ;
    inv02 ix64661 (.Y (nx64662), .A (nx65302)) ;
    inv02 ix64663 (.Y (nx64664), .A (nx65302)) ;
    inv02 ix64665 (.Y (nx64666), .A (nx65302)) ;
    inv02 ix64667 (.Y (nx64668), .A (nx65302)) ;
    inv02 ix64669 (.Y (nx64670), .A (nx65304)) ;
    inv02 ix64671 (.Y (nx64672), .A (nx65304)) ;
    inv02 ix64673 (.Y (nx64674), .A (nx65304)) ;
    inv02 ix64675 (.Y (nx64676), .A (nx65304)) ;
    inv02 ix64677 (.Y (nx64678), .A (nx238)) ;
    inv02 ix64679 (.Y (nx64680), .A (nx65294)) ;
    inv02 ix64681 (.Y (nx64682), .A (nx65294)) ;
    inv02 ix64683 (.Y (nx64684), .A (nx65294)) ;
    inv02 ix64685 (.Y (nx64686), .A (nx65294)) ;
    inv02 ix64687 (.Y (nx64688), .A (nx65294)) ;
    inv02 ix64689 (.Y (nx64690), .A (nx65294)) ;
    inv02 ix64691 (.Y (nx64692), .A (nx65294)) ;
    inv02 ix64693 (.Y (nx64694), .A (nx65296)) ;
    inv02 ix64695 (.Y (nx64696), .A (nx65296)) ;
    inv02 ix64697 (.Y (nx64698), .A (nx65296)) ;
    inv02 ix64699 (.Y (nx64700), .A (nx65296)) ;
    inv02 ix64701 (.Y (nx64702), .A (nx65296)) ;
    inv02 ix64703 (.Y (nx64704), .A (nx65296)) ;
    inv02 ix64705 (.Y (nx64706), .A (nx65296)) ;
    inv02 ix64707 (.Y (nx64708), .A (nx65298)) ;
    inv02 ix64709 (.Y (nx64710), .A (nx65298)) ;
    inv02 ix64711 (.Y (nx64712), .A (nx65298)) ;
    inv02 ix64713 (.Y (nx64714), .A (nx65298)) ;
    inv02 ix64715 (.Y (nx64716), .A (nx200)) ;
    inv02 ix64717 (.Y (nx64718), .A (nx65282)) ;
    inv02 ix64719 (.Y (nx64720), .A (nx65282)) ;
    inv02 ix64721 (.Y (nx64722), .A (nx65282)) ;
    inv02 ix64723 (.Y (nx64724), .A (nx65282)) ;
    inv02 ix64725 (.Y (nx64726), .A (nx65282)) ;
    inv02 ix64727 (.Y (nx64728), .A (nx65282)) ;
    inv02 ix64729 (.Y (nx64730), .A (nx65282)) ;
    inv02 ix64731 (.Y (nx64732), .A (nx65284)) ;
    inv02 ix64733 (.Y (nx64734), .A (nx65284)) ;
    inv02 ix64735 (.Y (nx64736), .A (nx65284)) ;
    inv02 ix64737 (.Y (nx64738), .A (nx65284)) ;
    inv02 ix64739 (.Y (nx64740), .A (nx65284)) ;
    inv02 ix64741 (.Y (nx64742), .A (nx65284)) ;
    inv02 ix64743 (.Y (nx64744), .A (nx65284)) ;
    inv02 ix64745 (.Y (nx64746), .A (nx65286)) ;
    inv02 ix64747 (.Y (nx64748), .A (nx65286)) ;
    inv02 ix64749 (.Y (nx64750), .A (nx65286)) ;
    inv02 ix64751 (.Y (nx64752), .A (nx65286)) ;
    inv02 ix64753 (.Y (nx64754), .A (nx218)) ;
    inv02 ix64755 (.Y (nx64756), .A (nx65288)) ;
    inv02 ix64757 (.Y (nx64758), .A (nx65288)) ;
    inv02 ix64759 (.Y (nx64760), .A (nx65288)) ;
    inv02 ix64761 (.Y (nx64762), .A (nx65288)) ;
    inv02 ix64763 (.Y (nx64764), .A (nx65288)) ;
    inv02 ix64765 (.Y (nx64766), .A (nx65288)) ;
    inv02 ix64767 (.Y (nx64768), .A (nx65288)) ;
    inv02 ix64769 (.Y (nx64770), .A (nx65290)) ;
    inv02 ix64771 (.Y (nx64772), .A (nx65290)) ;
    inv02 ix64773 (.Y (nx64774), .A (nx65290)) ;
    inv02 ix64775 (.Y (nx64776), .A (nx65290)) ;
    inv02 ix64777 (.Y (nx64778), .A (nx65290)) ;
    inv02 ix64779 (.Y (nx64780), .A (nx65290)) ;
    inv02 ix64781 (.Y (nx64782), .A (nx65290)) ;
    inv02 ix64783 (.Y (nx64784), .A (nx65292)) ;
    inv02 ix64785 (.Y (nx64786), .A (nx65292)) ;
    inv02 ix64787 (.Y (nx64788), .A (nx65292)) ;
    inv02 ix64789 (.Y (nx64790), .A (nx65292)) ;
    inv02 ix64791 (.Y (nx64792), .A (nx172)) ;
    inv02 ix64793 (.Y (nx64794), .A (nx65276)) ;
    inv02 ix64795 (.Y (nx64796), .A (nx65276)) ;
    inv02 ix64797 (.Y (nx64798), .A (nx65276)) ;
    inv02 ix64799 (.Y (nx64800), .A (nx65276)) ;
    inv02 ix64801 (.Y (nx64802), .A (nx65276)) ;
    inv02 ix64803 (.Y (nx64804), .A (nx65276)) ;
    inv02 ix64805 (.Y (nx64806), .A (nx65276)) ;
    inv02 ix64807 (.Y (nx64808), .A (nx65278)) ;
    inv02 ix64809 (.Y (nx64810), .A (nx65278)) ;
    inv02 ix64811 (.Y (nx64812), .A (nx65278)) ;
    inv02 ix64813 (.Y (nx64814), .A (nx65278)) ;
    inv02 ix64815 (.Y (nx64816), .A (nx65278)) ;
    inv02 ix64817 (.Y (nx64818), .A (nx65278)) ;
    inv02 ix64819 (.Y (nx64820), .A (nx65278)) ;
    inv02 ix64821 (.Y (nx64822), .A (nx65280)) ;
    inv02 ix64823 (.Y (nx64824), .A (nx65280)) ;
    inv02 ix64825 (.Y (nx64826), .A (nx65280)) ;
    inv02 ix64827 (.Y (nx64828), .A (nx65280)) ;
    inv02 ix64829 (.Y (nx64830), .A (nx154)) ;
    inv02 ix64831 (.Y (nx64832), .A (nx65270)) ;
    inv02 ix64833 (.Y (nx64834), .A (nx65270)) ;
    inv02 ix64835 (.Y (nx64836), .A (nx65270)) ;
    inv02 ix64837 (.Y (nx64838), .A (nx65270)) ;
    inv02 ix64839 (.Y (nx64840), .A (nx65270)) ;
    inv02 ix64841 (.Y (nx64842), .A (nx65270)) ;
    inv02 ix64843 (.Y (nx64844), .A (nx65270)) ;
    inv02 ix64845 (.Y (nx64846), .A (nx65272)) ;
    inv02 ix64847 (.Y (nx64848), .A (nx65272)) ;
    inv02 ix64849 (.Y (nx64850), .A (nx65272)) ;
    inv02 ix64851 (.Y (nx64852), .A (nx65272)) ;
    inv02 ix64853 (.Y (nx64854), .A (nx65272)) ;
    inv02 ix64855 (.Y (nx64856), .A (nx65272)) ;
    inv02 ix64857 (.Y (nx64858), .A (nx65272)) ;
    inv02 ix64859 (.Y (nx64860), .A (nx65274)) ;
    inv02 ix64861 (.Y (nx64862), .A (nx65274)) ;
    inv02 ix64863 (.Y (nx64864), .A (nx65274)) ;
    inv02 ix64865 (.Y (nx64866), .A (nx65274)) ;
    inv02 ix64867 (.Y (nx64868), .A (nx116)) ;
    inv02 ix64869 (.Y (nx64870), .A (nx65258)) ;
    inv02 ix64871 (.Y (nx64872), .A (nx65258)) ;
    inv02 ix64873 (.Y (nx64874), .A (nx65258)) ;
    inv02 ix64875 (.Y (nx64876), .A (nx65258)) ;
    inv02 ix64877 (.Y (nx64878), .A (nx65258)) ;
    inv02 ix64879 (.Y (nx64880), .A (nx65258)) ;
    inv02 ix64881 (.Y (nx64882), .A (nx65258)) ;
    inv02 ix64883 (.Y (nx64884), .A (nx65260)) ;
    inv02 ix64885 (.Y (nx64886), .A (nx65260)) ;
    inv02 ix64887 (.Y (nx64888), .A (nx65260)) ;
    inv02 ix64889 (.Y (nx64890), .A (nx65260)) ;
    inv02 ix64891 (.Y (nx64892), .A (nx65260)) ;
    inv02 ix64893 (.Y (nx64894), .A (nx65260)) ;
    inv02 ix64895 (.Y (nx64896), .A (nx65260)) ;
    inv02 ix64897 (.Y (nx64898), .A (nx65262)) ;
    inv02 ix64899 (.Y (nx64900), .A (nx65262)) ;
    inv02 ix64901 (.Y (nx64902), .A (nx65262)) ;
    inv02 ix64903 (.Y (nx64904), .A (nx65262)) ;
    inv02 ix64905 (.Y (nx64906), .A (nx134)) ;
    inv02 ix64907 (.Y (nx64908), .A (nx65264)) ;
    inv02 ix64909 (.Y (nx64910), .A (nx65264)) ;
    inv02 ix64911 (.Y (nx64912), .A (nx65264)) ;
    inv02 ix64913 (.Y (nx64914), .A (nx65264)) ;
    inv02 ix64915 (.Y (nx64916), .A (nx65264)) ;
    inv02 ix64917 (.Y (nx64918), .A (nx65264)) ;
    inv02 ix64919 (.Y (nx64920), .A (nx65264)) ;
    inv02 ix64921 (.Y (nx64922), .A (nx65266)) ;
    inv02 ix64923 (.Y (nx64924), .A (nx65266)) ;
    inv02 ix64925 (.Y (nx64926), .A (nx65266)) ;
    inv02 ix64927 (.Y (nx64928), .A (nx65266)) ;
    inv02 ix64929 (.Y (nx64930), .A (nx65266)) ;
    inv02 ix64931 (.Y (nx64932), .A (nx65266)) ;
    inv02 ix64933 (.Y (nx64934), .A (nx65266)) ;
    inv02 ix64935 (.Y (nx64936), .A (nx65268)) ;
    inv02 ix64937 (.Y (nx64938), .A (nx65268)) ;
    inv02 ix64939 (.Y (nx64940), .A (nx65268)) ;
    inv02 ix64941 (.Y (nx64942), .A (nx65268)) ;
    inv02 ix64943 (.Y (nx64944), .A (nx90)) ;
    inv02 ix64945 (.Y (nx64946), .A (nx65252)) ;
    inv02 ix64947 (.Y (nx64948), .A (nx65252)) ;
    inv02 ix64949 (.Y (nx64950), .A (nx65252)) ;
    inv02 ix64951 (.Y (nx64952), .A (nx65252)) ;
    inv02 ix64953 (.Y (nx64954), .A (nx65252)) ;
    inv02 ix64955 (.Y (nx64956), .A (nx65252)) ;
    inv02 ix64957 (.Y (nx64958), .A (nx65252)) ;
    inv02 ix64959 (.Y (nx64960), .A (nx65254)) ;
    inv02 ix64961 (.Y (nx64962), .A (nx65254)) ;
    inv02 ix64963 (.Y (nx64964), .A (nx65254)) ;
    inv02 ix64965 (.Y (nx64966), .A (nx65254)) ;
    inv02 ix64967 (.Y (nx64968), .A (nx65254)) ;
    inv02 ix64969 (.Y (nx64970), .A (nx65254)) ;
    inv02 ix64971 (.Y (nx64972), .A (nx65254)) ;
    inv02 ix64973 (.Y (nx64974), .A (nx65256)) ;
    inv02 ix64975 (.Y (nx64976), .A (nx65256)) ;
    inv02 ix64977 (.Y (nx64978), .A (nx65256)) ;
    inv02 ix64979 (.Y (nx64980), .A (nx65256)) ;
    inv02 ix64981 (.Y (nx64982), .A (nx70)) ;
    inv02 ix64983 (.Y (nx64984), .A (nx65246)) ;
    inv02 ix64985 (.Y (nx64986), .A (nx65246)) ;
    inv02 ix64987 (.Y (nx64988), .A (nx65246)) ;
    inv02 ix64989 (.Y (nx64990), .A (nx65246)) ;
    inv02 ix64991 (.Y (nx64992), .A (nx65246)) ;
    inv02 ix64993 (.Y (nx64994), .A (nx65246)) ;
    inv02 ix64995 (.Y (nx64996), .A (nx65246)) ;
    inv02 ix64997 (.Y (nx64998), .A (nx65248)) ;
    inv02 ix64999 (.Y (nx65000), .A (nx65248)) ;
    inv02 ix65001 (.Y (nx65002), .A (nx65248)) ;
    inv02 ix65003 (.Y (nx65004), .A (nx65248)) ;
    inv02 ix65005 (.Y (nx65006), .A (nx65248)) ;
    inv02 ix65007 (.Y (nx65008), .A (nx65248)) ;
    inv02 ix65009 (.Y (nx65010), .A (nx65248)) ;
    inv02 ix65011 (.Y (nx65012), .A (nx65250)) ;
    inv02 ix65013 (.Y (nx65014), .A (nx65250)) ;
    inv02 ix65015 (.Y (nx65016), .A (nx65250)) ;
    inv02 ix65017 (.Y (nx65018), .A (nx65250)) ;
    inv02 ix65019 (.Y (nx65020), .A (nx24)) ;
    inv02 ix65021 (.Y (nx65022), .A (nx65234)) ;
    inv02 ix65023 (.Y (nx65024), .A (nx65234)) ;
    inv02 ix65025 (.Y (nx65026), .A (nx65234)) ;
    inv02 ix65027 (.Y (nx65028), .A (nx65234)) ;
    inv02 ix65029 (.Y (nx65030), .A (nx65234)) ;
    inv02 ix65031 (.Y (nx65032), .A (nx65234)) ;
    inv02 ix65033 (.Y (nx65034), .A (nx65234)) ;
    inv02 ix65035 (.Y (nx65036), .A (nx65236)) ;
    inv02 ix65037 (.Y (nx65038), .A (nx65236)) ;
    inv02 ix65039 (.Y (nx65040), .A (nx65236)) ;
    inv02 ix65041 (.Y (nx65042), .A (nx65236)) ;
    inv02 ix65043 (.Y (nx65044), .A (nx65236)) ;
    inv02 ix65045 (.Y (nx65046), .A (nx65236)) ;
    inv02 ix65047 (.Y (nx65048), .A (nx65236)) ;
    inv02 ix65049 (.Y (nx65050), .A (nx65238)) ;
    inv02 ix65051 (.Y (nx65052), .A (nx65238)) ;
    inv02 ix65053 (.Y (nx65054), .A (nx65238)) ;
    inv02 ix65055 (.Y (nx65056), .A (nx65238)) ;
    inv02 ix65057 (.Y (nx65058), .A (nx46)) ;
    inv02 ix65059 (.Y (nx65060), .A (nx65240)) ;
    inv02 ix65061 (.Y (nx65062), .A (nx65240)) ;
    inv02 ix65063 (.Y (nx65064), .A (nx65240)) ;
    inv02 ix65065 (.Y (nx65066), .A (nx65240)) ;
    inv02 ix65067 (.Y (nx65068), .A (nx65240)) ;
    inv02 ix65069 (.Y (nx65070), .A (nx65240)) ;
    inv02 ix65071 (.Y (nx65072), .A (nx65240)) ;
    inv02 ix65073 (.Y (nx65074), .A (nx65242)) ;
    inv02 ix65075 (.Y (nx65076), .A (nx65242)) ;
    inv02 ix65077 (.Y (nx65078), .A (nx65242)) ;
    inv02 ix65079 (.Y (nx65080), .A (nx65242)) ;
    inv02 ix65081 (.Y (nx65082), .A (nx65242)) ;
    inv02 ix65083 (.Y (nx65084), .A (nx65242)) ;
    inv02 ix65085 (.Y (nx65086), .A (nx65242)) ;
    inv02 ix65087 (.Y (nx65088), .A (nx65244)) ;
    inv02 ix65089 (.Y (nx65090), .A (nx65244)) ;
    inv02 ix65091 (.Y (nx65092), .A (nx65244)) ;
    inv02 ix65093 (.Y (nx65094), .A (nx65244)) ;
    inv02 ix65095 (.Y (nx65096), .A (nx4498)) ;
    inv02 ix65097 (.Y (nx65098), .A (nx4498)) ;
    inv02 ix65099 (.Y (nx65100), .A (nx4206)) ;
    inv02 ix65101 (.Y (nx65102), .A (nx4206)) ;
    inv02 ix65103 (.Y (nx65104), .A (nx3912)) ;
    inv02 ix65105 (.Y (nx65106), .A (nx3912)) ;
    inv02 ix65107 (.Y (nx65108), .A (nx3620)) ;
    inv02 ix65109 (.Y (nx65110), .A (nx3620)) ;
    inv02 ix65111 (.Y (nx65112), .A (nx3318)) ;
    inv02 ix65113 (.Y (nx65114), .A (nx3318)) ;
    inv02 ix65115 (.Y (nx65116), .A (nx3026)) ;
    inv02 ix65117 (.Y (nx65118), .A (nx3026)) ;
    inv02 ix65119 (.Y (nx65120), .A (nx2732)) ;
    inv02 ix65121 (.Y (nx65122), .A (nx2732)) ;
    inv02 ix65123 (.Y (nx65124), .A (nx2440)) ;
    inv02 ix65125 (.Y (nx65126), .A (nx2440)) ;
    inv02 ix65127 (.Y (nx65128), .A (nx2142)) ;
    inv02 ix65129 (.Y (nx65130), .A (nx2142)) ;
    buf02 ix65131 (.Y (nx65132), .A (nx54994)) ;
    buf02 ix65133 (.Y (nx65134), .A (nx54994)) ;
    inv01 ix65135 (.Y (nx65136), .A (nx54996)) ;
    inv02 ix65137 (.Y (nx65138), .A (nx65136)) ;
    inv02 ix65139 (.Y (nx65140), .A (nx65136)) ;
    inv02 ix65141 (.Y (nx65142), .A (nx65136)) ;
    inv02 ix65143 (.Y (nx65144), .A (nx65136)) ;
    buf02 ix65145 (.Y (nx65146), .A (nx55001)) ;
    buf02 ix65147 (.Y (nx65148), .A (nx55001)) ;
    buf02 ix65149 (.Y (nx65150), .A (nx55008)) ;
    buf02 ix65151 (.Y (nx65152), .A (nx55008)) ;
    buf02 ix65153 (.Y (nx65154), .A (nx55013)) ;
    buf02 ix65155 (.Y (nx65156), .A (nx55013)) ;
    buf02 ix65157 (.Y (nx65158), .A (nx55020)) ;
    buf02 ix65159 (.Y (nx65160), .A (nx55020)) ;
    buf02 ix65161 (.Y (nx65162), .A (nx55025)) ;
    buf02 ix65163 (.Y (nx65164), .A (nx55025)) ;
    buf02 ix65165 (.Y (nx65166), .A (nx55032)) ;
    buf02 ix65167 (.Y (nx65168), .A (nx55032)) ;
    buf02 ix65169 (.Y (nx65170), .A (nx55037)) ;
    buf02 ix65171 (.Y (nx65172), .A (nx55037)) ;
    buf02 ix65173 (.Y (nx65174), .A (nx55045)) ;
    buf02 ix65175 (.Y (nx65176), .A (nx55045)) ;
    buf02 ix65177 (.Y (nx65178), .A (nx55050)) ;
    buf02 ix65179 (.Y (nx65180), .A (nx55050)) ;
    buf02 ix65181 (.Y (nx65182), .A (nx55057)) ;
    buf02 ix65183 (.Y (nx65184), .A (nx55057)) ;
    buf02 ix65185 (.Y (nx65186), .A (nx55062)) ;
    buf02 ix65187 (.Y (nx65188), .A (nx55062)) ;
    buf02 ix65189 (.Y (nx65190), .A (nx55069)) ;
    buf02 ix65191 (.Y (nx65192), .A (nx55069)) ;
    buf02 ix65193 (.Y (nx65194), .A (nx55074)) ;
    buf02 ix65195 (.Y (nx65196), .A (nx55074)) ;
    buf02 ix65197 (.Y (nx65198), .A (nx55081)) ;
    buf02 ix65199 (.Y (nx65200), .A (nx55081)) ;
    buf02 ix65201 (.Y (nx65202), .A (nx55086)) ;
    buf02 ix65203 (.Y (nx65204), .A (nx55086)) ;
    inv02 ix65205 (.Y (nx65206), .A (nx1554)) ;
    inv02 ix65207 (.Y (nx65208), .A (nx1554)) ;
    inv02 ix65209 (.Y (nx65210), .A (nx1262)) ;
    inv02 ix65211 (.Y (nx65212), .A (nx1262)) ;
    inv02 ix65213 (.Y (nx65214), .A (nx962)) ;
    inv02 ix65215 (.Y (nx65216), .A (nx962)) ;
    inv02 ix65217 (.Y (nx65218), .A (nx668)) ;
    inv02 ix65219 (.Y (nx65220), .A (nx668)) ;
    inv02 ix65221 (.Y (nx65222), .A (nx370)) ;
    inv02 ix65223 (.Y (nx65224), .A (nx370)) ;
    inv02 ix65225 (.Y (nx65226), .A (nx10)) ;
    inv02 ix65227 (.Y (nx65228), .A (nx10)) ;
    inv02 ix65233 (.Y (nx65234), .A (nx65020)) ;
    inv02 ix65235 (.Y (nx65236), .A (nx65020)) ;
    inv02 ix65237 (.Y (nx65238), .A (nx65020)) ;
    inv02 ix65239 (.Y (nx65240), .A (nx65058)) ;
    inv02 ix65241 (.Y (nx65242), .A (nx65058)) ;
    inv02 ix65243 (.Y (nx65244), .A (nx65058)) ;
    inv02 ix65245 (.Y (nx65246), .A (nx64982)) ;
    inv02 ix65247 (.Y (nx65248), .A (nx64982)) ;
    inv02 ix65249 (.Y (nx65250), .A (nx64982)) ;
    inv02 ix65251 (.Y (nx65252), .A (nx64944)) ;
    inv02 ix65253 (.Y (nx65254), .A (nx64944)) ;
    inv02 ix65255 (.Y (nx65256), .A (nx64944)) ;
    inv02 ix65257 (.Y (nx65258), .A (nx64868)) ;
    inv02 ix65259 (.Y (nx65260), .A (nx64868)) ;
    inv02 ix65261 (.Y (nx65262), .A (nx64868)) ;
    inv02 ix65263 (.Y (nx65264), .A (nx64906)) ;
    inv02 ix65265 (.Y (nx65266), .A (nx64906)) ;
    inv02 ix65267 (.Y (nx65268), .A (nx64906)) ;
    inv02 ix65269 (.Y (nx65270), .A (nx64830)) ;
    inv02 ix65271 (.Y (nx65272), .A (nx64830)) ;
    inv02 ix65273 (.Y (nx65274), .A (nx64830)) ;
    inv02 ix65275 (.Y (nx65276), .A (nx64792)) ;
    inv02 ix65277 (.Y (nx65278), .A (nx64792)) ;
    inv02 ix65279 (.Y (nx65280), .A (nx64792)) ;
    inv02 ix65281 (.Y (nx65282), .A (nx64716)) ;
    inv02 ix65283 (.Y (nx65284), .A (nx64716)) ;
    inv02 ix65285 (.Y (nx65286), .A (nx64716)) ;
    inv02 ix65287 (.Y (nx65288), .A (nx64754)) ;
    inv02 ix65289 (.Y (nx65290), .A (nx64754)) ;
    inv02 ix65291 (.Y (nx65292), .A (nx64754)) ;
    inv02 ix65293 (.Y (nx65294), .A (nx64678)) ;
    inv02 ix65295 (.Y (nx65296), .A (nx64678)) ;
    inv02 ix65297 (.Y (nx65298), .A (nx64678)) ;
    inv02 ix65299 (.Y (nx65300), .A (nx64640)) ;
    inv02 ix65301 (.Y (nx65302), .A (nx64640)) ;
    inv02 ix65303 (.Y (nx65304), .A (nx64640)) ;
    inv02 ix65305 (.Y (nx65306), .A (nx64564)) ;
    inv02 ix65307 (.Y (nx65308), .A (nx64564)) ;
    inv02 ix65309 (.Y (nx65310), .A (nx64564)) ;
    inv02 ix65311 (.Y (nx65312), .A (nx64602)) ;
    inv02 ix65313 (.Y (nx65314), .A (nx64602)) ;
    inv02 ix65315 (.Y (nx65316), .A (nx64602)) ;
    inv02 ix65317 (.Y (nx65318), .A (nx64526)) ;
    inv02 ix65319 (.Y (nx65320), .A (nx64526)) ;
    inv02 ix65321 (.Y (nx65322), .A (nx64526)) ;
    inv02 ix65323 (.Y (nx65324), .A (nx54129)) ;
    inv02 ix65325 (.Y (nx65326), .A (nx54129)) ;
    inv02 ix65327 (.Y (nx65328), .A (nx54129)) ;
    inv02 ix65329 (.Y (nx65330), .A (nx318)) ;
    inv02 ix65331 (.Y (nx65332), .A (nx280)) ;
    inv02 ix65333 (.Y (nx65334), .A (nx298)) ;
    inv02 ix65335 (.Y (nx65336), .A (nx256)) ;
    inv02 ix65337 (.Y (nx65338), .A (nx238)) ;
    inv02 ix65339 (.Y (nx65340), .A (nx200)) ;
    inv02 ix65341 (.Y (nx65342), .A (nx218)) ;
    inv02 ix65343 (.Y (nx65344), .A (nx172)) ;
    inv02 ix65345 (.Y (nx65346), .A (nx154)) ;
    inv02 ix65347 (.Y (nx65348), .A (nx116)) ;
    inv02 ix65349 (.Y (nx65350), .A (nx134)) ;
    inv02 ix65351 (.Y (nx65352), .A (nx90)) ;
    inv02 ix65353 (.Y (nx65354), .A (nx70)) ;
    inv02 ix65355 (.Y (nx65356), .A (nx24)) ;
    inv02 ix65357 (.Y (nx65358), .A (nx46)) ;
    and03 ix4769 (.Y (nx4768), .A0 (nx66120), .A1 (nx65370), .A2 (nx66056)) ;
    and03 ix4753 (.Y (nx4752), .A0 (nx66120), .A1 (nx65370), .A2 (nx66060)) ;
    nor02ii ix54136 (.Y (nx54135), .A0 (nx65444), .A1 (address[0])) ;
    and03 ix4719 (.Y (nx4718), .A0 (nx66120), .A1 (nx65370), .A2 (nx66064)) ;
    and03 ix4735 (.Y (nx4734), .A0 (nx66120), .A1 (nx65370), .A2 (nx66068)) ;
    nor02ii ix54157 (.Y (nx54156), .A0 (address[0]), .A1 (nx65446)) ;
    and03 ix4699 (.Y (nx4698), .A0 (nx66120), .A1 (nx65370), .A2 (nx66072)) ;
    nor02ii ix54170 (.Y (nx54169), .A0 (address[3]), .A1 (address[2])) ;
    and03 ix4683 (.Y (nx4682), .A0 (nx66120), .A1 (nx65372), .A2 (nx66076)) ;
    and03 ix4649 (.Y (nx4648), .A0 (nx66122), .A1 (nx65372), .A2 (nx66080)) ;
    and03 ix4665 (.Y (nx4664), .A0 (nx66122), .A1 (nx65372), .A2 (nx66084)) ;
    and03 ix4627 (.Y (nx4626), .A0 (nx66122), .A1 (nx65372), .A2 (nx66088)) ;
    nor02ii ix54207 (.Y (nx54206), .A0 (address[2]), .A1 (address[3])) ;
    and03 ix4611 (.Y (nx4610), .A0 (nx66122), .A1 (nx65372), .A2 (nx66092)) ;
    and03 ix4577 (.Y (nx4576), .A0 (nx66122), .A1 (nx65372), .A2 (nx66096)) ;
    and03 ix4593 (.Y (nx4592), .A0 (nx66122), .A1 (nx65372), .A2 (nx66100)) ;
    and03 ix4557 (.Y (nx4556), .A0 (nx66122), .A1 (nx65374), .A2 (nx66104)) ;
    and03 ix4541 (.Y (nx4540), .A0 (nx65098), .A1 (nx65374), .A2 (nx66108)) ;
    and03 ix4507 (.Y (nx4506), .A0 (nx65098), .A1 (nx65374), .A2 (nx66112)) ;
    and03 ix4523 (.Y (nx4522), .A0 (nx65098), .A1 (nx65374), .A2 (nx66116)) ;
    and03 ix4477 (.Y (nx4476), .A0 (nx66124), .A1 (nx65374), .A2 (nx66056)) ;
    nor02ii ix54283 (.Y (nx54282), .A0 (address[4]), .A1 (nx65440)) ;
    and03 ix4461 (.Y (nx4460), .A0 (nx66124), .A1 (nx65374), .A2 (nx66060)) ;
    and03 ix4427 (.Y (nx4426), .A0 (nx66124), .A1 (nx65374), .A2 (nx66064)) ;
    and03 ix4443 (.Y (nx4442), .A0 (nx66124), .A1 (nx65376), .A2 (nx66068)) ;
    and03 ix4407 (.Y (nx4406), .A0 (nx66124), .A1 (nx65376), .A2 (nx66072)) ;
    and03 ix4391 (.Y (nx4390), .A0 (nx66124), .A1 (nx65376), .A2 (nx66076)) ;
    and03 ix4357 (.Y (nx4356), .A0 (nx66126), .A1 (nx65376), .A2 (nx66080)) ;
    and03 ix4373 (.Y (nx4372), .A0 (nx66126), .A1 (nx65376), .A2 (nx66084)) ;
    and03 ix4335 (.Y (nx4334), .A0 (nx66126), .A1 (nx65376), .A2 (nx66088)) ;
    and03 ix4319 (.Y (nx4318), .A0 (nx66126), .A1 (nx65376), .A2 (nx66092)) ;
    and03 ix4285 (.Y (nx4284), .A0 (nx66126), .A1 (nx65378), .A2 (nx66096)) ;
    and03 ix4301 (.Y (nx4300), .A0 (nx66126), .A1 (nx65378), .A2 (nx66100)) ;
    and03 ix4265 (.Y (nx4264), .A0 (nx66126), .A1 (nx65378), .A2 (nx66104)) ;
    and03 ix4249 (.Y (nx4248), .A0 (nx65102), .A1 (nx65378), .A2 (nx66108)) ;
    and03 ix4215 (.Y (nx4214), .A0 (nx65102), .A1 (nx65378), .A2 (nx66112)) ;
    and03 ix4231 (.Y (nx4230), .A0 (nx65102), .A1 (nx65378), .A2 (nx66116)) ;
    and03 ix4183 (.Y (nx4182), .A0 (nx66128), .A1 (nx65378), .A2 (nx66056)) ;
    nor02ii ix54374 (.Y (nx54373), .A0 (nx65442), .A1 (address[4])) ;
    and03 ix4167 (.Y (nx4166), .A0 (nx66128), .A1 (nx65380), .A2 (nx66060)) ;
    and03 ix4133 (.Y (nx4132), .A0 (nx66128), .A1 (nx65380), .A2 (nx66064)) ;
    and03 ix4149 (.Y (nx4148), .A0 (nx66128), .A1 (nx65380), .A2 (nx66068)) ;
    and03 ix4113 (.Y (nx4112), .A0 (nx66128), .A1 (nx65380), .A2 (nx66072)) ;
    and03 ix4097 (.Y (nx4096), .A0 (nx66128), .A1 (nx65380), .A2 (nx66076)) ;
    and03 ix4063 (.Y (nx4062), .A0 (nx66130), .A1 (nx65380), .A2 (nx66080)) ;
    and03 ix4079 (.Y (nx4078), .A0 (nx66130), .A1 (nx65380), .A2 (nx66084)) ;
    and03 ix4041 (.Y (nx4040), .A0 (nx66130), .A1 (nx65382), .A2 (nx66088)) ;
    and03 ix4025 (.Y (nx4024), .A0 (nx66130), .A1 (nx65382), .A2 (nx66092)) ;
    and03 ix3991 (.Y (nx3990), .A0 (nx66130), .A1 (nx65382), .A2 (nx66096)) ;
    and03 ix4007 (.Y (nx4006), .A0 (nx66130), .A1 (nx65382), .A2 (nx66100)) ;
    and03 ix3971 (.Y (nx3970), .A0 (nx66130), .A1 (nx65382), .A2 (nx66104)) ;
    and03 ix3955 (.Y (nx3954), .A0 (nx65106), .A1 (nx65382), .A2 (nx66108)) ;
    and03 ix3921 (.Y (nx3920), .A0 (nx65106), .A1 (nx65382), .A2 (nx66112)) ;
    and03 ix3937 (.Y (nx3936), .A0 (nx65106), .A1 (nx65384), .A2 (nx66116)) ;
    and03 ix3891 (.Y (nx3890), .A0 (nx66132), .A1 (nx65384), .A2 (nx66056)) ;
    and03 ix3875 (.Y (nx3874), .A0 (nx66132), .A1 (nx65384), .A2 (nx66060)) ;
    and03 ix3841 (.Y (nx3840), .A0 (nx66132), .A1 (nx65384), .A2 (nx66064)) ;
    and03 ix3857 (.Y (nx3856), .A0 (nx66132), .A1 (nx65384), .A2 (nx66068)) ;
    and03 ix3821 (.Y (nx3820), .A0 (nx66132), .A1 (nx65384), .A2 (nx66072)) ;
    and03 ix3805 (.Y (nx3804), .A0 (nx66132), .A1 (nx65384), .A2 (nx66076)) ;
    and03 ix3771 (.Y (nx3770), .A0 (nx66134), .A1 (nx65386), .A2 (nx66080)) ;
    and03 ix3787 (.Y (nx3786), .A0 (nx66134), .A1 (nx65386), .A2 (nx66084)) ;
    and03 ix3749 (.Y (nx3748), .A0 (nx66134), .A1 (nx65386), .A2 (nx66088)) ;
    and03 ix3733 (.Y (nx3732), .A0 (nx66134), .A1 (nx65386), .A2 (nx66092)) ;
    and03 ix3699 (.Y (nx3698), .A0 (nx66134), .A1 (nx65386), .A2 (nx66096)) ;
    and03 ix3715 (.Y (nx3714), .A0 (nx66134), .A1 (nx65386), .A2 (nx66100)) ;
    and03 ix3679 (.Y (nx3678), .A0 (nx66134), .A1 (nx65386), .A2 (nx66104)) ;
    and03 ix3663 (.Y (nx3662), .A0 (nx65110), .A1 (nx65388), .A2 (nx66108)) ;
    and03 ix3629 (.Y (nx3628), .A0 (nx65110), .A1 (nx65388), .A2 (nx66112)) ;
    and03 ix3645 (.Y (nx3644), .A0 (nx65110), .A1 (nx65388), .A2 (nx66116)) ;
    and03 ix3589 (.Y (nx3588), .A0 (nx66136), .A1 (nx65388), .A2 (nx66058)) ;
    nor02ii ix54555 (.Y (nx54554), .A0 (address[7]), .A1 (address[6])) ;
    and03 ix3573 (.Y (nx3572), .A0 (nx66136), .A1 (nx65388), .A2 (nx66062)) ;
    and03 ix3539 (.Y (nx3538), .A0 (nx66136), .A1 (nx65388), .A2 (nx66066)) ;
    and03 ix3555 (.Y (nx3554), .A0 (nx66136), .A1 (nx65388), .A2 (nx66070)) ;
    and03 ix3519 (.Y (nx3518), .A0 (nx66136), .A1 (nx65390), .A2 (nx66074)) ;
    and03 ix3503 (.Y (nx3502), .A0 (nx66136), .A1 (nx65390), .A2 (nx66078)) ;
    and03 ix3469 (.Y (nx3468), .A0 (nx66138), .A1 (nx65390), .A2 (nx66082)) ;
    and03 ix3485 (.Y (nx3484), .A0 (nx66138), .A1 (nx65390), .A2 (nx66086)) ;
    and03 ix3447 (.Y (nx3446), .A0 (nx66138), .A1 (nx65390), .A2 (nx66090)) ;
    and03 ix3431 (.Y (nx3430), .A0 (nx66138), .A1 (nx65390), .A2 (nx66094)) ;
    and03 ix3397 (.Y (nx3396), .A0 (nx66138), .A1 (nx65390), .A2 (nx66098)) ;
    and03 ix3413 (.Y (nx3412), .A0 (nx66138), .A1 (nx65392), .A2 (nx66102)) ;
    and03 ix3377 (.Y (nx3376), .A0 (nx66138), .A1 (nx65392), .A2 (nx66106)) ;
    and03 ix3361 (.Y (nx3360), .A0 (nx65114), .A1 (nx65392), .A2 (nx66110)) ;
    and03 ix3327 (.Y (nx3326), .A0 (nx65114), .A1 (nx65392), .A2 (nx66114)) ;
    and03 ix3343 (.Y (nx3342), .A0 (nx65114), .A1 (nx65392), .A2 (nx66118)) ;
    and03 ix3297 (.Y (nx3296), .A0 (nx66140), .A1 (nx65392), .A2 (nx66058)) ;
    and03 ix3281 (.Y (nx3280), .A0 (nx66140), .A1 (nx65392), .A2 (nx66062)) ;
    and03 ix3247 (.Y (nx3246), .A0 (nx66140), .A1 (nx65394), .A2 (nx66066)) ;
    and03 ix3263 (.Y (nx3262), .A0 (nx66140), .A1 (nx65394), .A2 (nx66070)) ;
    and03 ix3227 (.Y (nx3226), .A0 (nx66140), .A1 (nx65394), .A2 (nx66074)) ;
    and03 ix3211 (.Y (nx3210), .A0 (nx66140), .A1 (nx65394), .A2 (nx66078)) ;
    and03 ix3177 (.Y (nx3176), .A0 (nx66142), .A1 (nx65394), .A2 (nx66082)) ;
    and03 ix3193 (.Y (nx3192), .A0 (nx66142), .A1 (nx65394), .A2 (nx66086)) ;
    and03 ix3155 (.Y (nx3154), .A0 (nx66142), .A1 (nx65394), .A2 (nx66090)) ;
    and03 ix3139 (.Y (nx3138), .A0 (nx66142), .A1 (nx65396), .A2 (nx66094)) ;
    and03 ix3105 (.Y (nx3104), .A0 (nx66142), .A1 (nx65396), .A2 (nx66098)) ;
    and03 ix3121 (.Y (nx3120), .A0 (nx66142), .A1 (nx65396), .A2 (nx66102)) ;
    and03 ix3085 (.Y (nx3084), .A0 (nx66142), .A1 (nx65396), .A2 (nx66106)) ;
    and03 ix3069 (.Y (nx3068), .A0 (nx65118), .A1 (nx65396), .A2 (nx66110)) ;
    and03 ix3035 (.Y (nx3034), .A0 (nx65118), .A1 (nx65396), .A2 (nx66114)) ;
    and03 ix3051 (.Y (nx3050), .A0 (nx65118), .A1 (nx65396), .A2 (nx66118)) ;
    and03 ix3003 (.Y (nx3002), .A0 (nx66144), .A1 (nx65398), .A2 (nx66058)) ;
    and03 ix2987 (.Y (nx2986), .A0 (nx66144), .A1 (nx65398), .A2 (nx66062)) ;
    and03 ix2953 (.Y (nx2952), .A0 (nx66144), .A1 (nx65398), .A2 (nx66066)) ;
    and03 ix2969 (.Y (nx2968), .A0 (nx66144), .A1 (nx65398), .A2 (nx66070)) ;
    and03 ix2933 (.Y (nx2932), .A0 (nx66144), .A1 (nx65398), .A2 (nx66074)) ;
    and03 ix2917 (.Y (nx2916), .A0 (nx66144), .A1 (nx65398), .A2 (nx66078)) ;
    and03 ix2883 (.Y (nx2882), .A0 (nx66146), .A1 (nx65398), .A2 (nx66082)) ;
    and03 ix2899 (.Y (nx2898), .A0 (nx66146), .A1 (nx65400), .A2 (nx66086)) ;
    and03 ix2861 (.Y (nx2860), .A0 (nx66146), .A1 (nx65400), .A2 (nx66090)) ;
    and03 ix2845 (.Y (nx2844), .A0 (nx66146), .A1 (nx65400), .A2 (nx66094)) ;
    and03 ix2811 (.Y (nx2810), .A0 (nx66146), .A1 (nx65400), .A2 (nx66098)) ;
    and03 ix2827 (.Y (nx2826), .A0 (nx66146), .A1 (nx65400), .A2 (nx66102)) ;
    and03 ix2791 (.Y (nx2790), .A0 (nx66146), .A1 (nx65400), .A2 (nx66106)) ;
    and03 ix2775 (.Y (nx2774), .A0 (nx65122), .A1 (nx65400), .A2 (nx66110)) ;
    and03 ix2741 (.Y (nx2740), .A0 (nx65122), .A1 (nx65402), .A2 (nx66114)) ;
    and03 ix2757 (.Y (nx2756), .A0 (nx65122), .A1 (nx65402), .A2 (nx66118)) ;
    and03 ix2711 (.Y (nx2710), .A0 (nx66148), .A1 (nx65402), .A2 (nx66058)) ;
    and03 ix2695 (.Y (nx2694), .A0 (nx66148), .A1 (nx65402), .A2 (nx66062)) ;
    and03 ix2661 (.Y (nx2660), .A0 (nx66148), .A1 (nx65402), .A2 (nx66066)) ;
    and03 ix2677 (.Y (nx2676), .A0 (nx66148), .A1 (nx65402), .A2 (nx66070)) ;
    and03 ix2641 (.Y (nx2640), .A0 (nx66148), .A1 (nx65402), .A2 (nx66074)) ;
    and03 ix2625 (.Y (nx2624), .A0 (nx66148), .A1 (nx65404), .A2 (nx66078)) ;
    and03 ix2591 (.Y (nx2590), .A0 (nx66150), .A1 (nx65404), .A2 (nx66082)) ;
    and03 ix2607 (.Y (nx2606), .A0 (nx66150), .A1 (nx65404), .A2 (nx66086)) ;
    and03 ix2569 (.Y (nx2568), .A0 (nx66150), .A1 (nx65404), .A2 (nx66090)) ;
    and03 ix2553 (.Y (nx2552), .A0 (nx66150), .A1 (nx65404), .A2 (nx66094)) ;
    and03 ix2519 (.Y (nx2518), .A0 (nx66150), .A1 (nx65404), .A2 (nx66098)) ;
    and03 ix2535 (.Y (nx2534), .A0 (nx66150), .A1 (nx65404), .A2 (nx66102)) ;
    and03 ix2499 (.Y (nx2498), .A0 (nx66150), .A1 (nx65406), .A2 (nx66106)) ;
    and03 ix2483 (.Y (nx2482), .A0 (nx65126), .A1 (nx65406), .A2 (nx66110)) ;
    and03 ix2449 (.Y (nx2448), .A0 (nx65126), .A1 (nx65406), .A2 (nx66114)) ;
    and03 ix2465 (.Y (nx2464), .A0 (nx65126), .A1 (nx65406), .A2 (nx66118)) ;
    and03 ix2413 (.Y (nx2412), .A0 (nx66152), .A1 (nx65406), .A2 (nx66058)) ;
    and03 ix2397 (.Y (nx2396), .A0 (nx66152), .A1 (nx65406), .A2 (nx66062)) ;
    and03 ix2363 (.Y (nx2362), .A0 (nx66152), .A1 (nx65406), .A2 (nx66066)) ;
    and03 ix2379 (.Y (nx2378), .A0 (nx66152), .A1 (nx65408), .A2 (nx66070)) ;
    and03 ix2343 (.Y (nx2342), .A0 (nx66152), .A1 (nx65408), .A2 (nx66074)) ;
    and03 ix2327 (.Y (nx2326), .A0 (nx66152), .A1 (nx65408), .A2 (nx66078)) ;
    and03 ix2293 (.Y (nx2292), .A0 (nx66154), .A1 (nx65408), .A2 (nx66082)) ;
    and03 ix2309 (.Y (nx2308), .A0 (nx66154), .A1 (nx65408), .A2 (nx66086)) ;
    and03 ix2271 (.Y (nx2270), .A0 (nx66154), .A1 (nx65408), .A2 (nx66090)) ;
    and03 ix2255 (.Y (nx2254), .A0 (nx66154), .A1 (nx65408), .A2 (nx66094)) ;
    and03 ix2221 (.Y (nx2220), .A0 (nx66154), .A1 (nx65410), .A2 (nx66098)) ;
    and03 ix2237 (.Y (nx2236), .A0 (nx66154), .A1 (nx65410), .A2 (nx66102)) ;
    and03 ix2201 (.Y (nx2200), .A0 (nx66154), .A1 (nx65410), .A2 (nx66106)) ;
    and03 ix2185 (.Y (nx2184), .A0 (nx65130), .A1 (nx65410), .A2 (nx66110)) ;
    and03 ix2151 (.Y (nx2150), .A0 (nx65130), .A1 (nx65410), .A2 (nx66114)) ;
    and03 ix2167 (.Y (nx2166), .A0 (nx65130), .A1 (nx65410), .A2 (nx66118)) ;
    and03 ix1825 (.Y (nx1824), .A0 (nx66156), .A1 (nx65410), .A2 (nx66058)) ;
    and03 ix1809 (.Y (nx1808), .A0 (nx66156), .A1 (nx65412), .A2 (nx66062)) ;
    and03 ix1775 (.Y (nx1774), .A0 (nx66156), .A1 (nx65412), .A2 (nx66066)) ;
    and03 ix1791 (.Y (nx1790), .A0 (nx66156), .A1 (nx65412), .A2 (nx66070)) ;
    and03 ix1755 (.Y (nx1754), .A0 (nx66156), .A1 (nx65412), .A2 (nx66074)) ;
    and03 ix1739 (.Y (nx1738), .A0 (nx66156), .A1 (nx65412), .A2 (nx66078)) ;
    and03 ix1705 (.Y (nx1704), .A0 (nx66158), .A1 (nx65412), .A2 (nx66082)) ;
    and03 ix1721 (.Y (nx1720), .A0 (nx66158), .A1 (nx65412), .A2 (nx66086)) ;
    and03 ix1683 (.Y (nx1682), .A0 (nx66158), .A1 (nx65414), .A2 (nx66090)) ;
    and03 ix1667 (.Y (nx1666), .A0 (nx66158), .A1 (nx65414), .A2 (nx66094)) ;
    and03 ix1633 (.Y (nx1632), .A0 (nx66158), .A1 (nx65414), .A2 (nx66098)) ;
    and03 ix1649 (.Y (nx1648), .A0 (nx66158), .A1 (nx65414), .A2 (nx66102)) ;
    and03 ix1613 (.Y (nx1612), .A0 (nx66158), .A1 (nx65414), .A2 (nx66106)) ;
    and03 ix1597 (.Y (nx1596), .A0 (nx65208), .A1 (nx65414), .A2 (nx66110)) ;
    and03 ix1563 (.Y (nx1562), .A0 (nx65208), .A1 (nx65414), .A2 (nx66114)) ;
    and03 ix1579 (.Y (nx1578), .A0 (nx65208), .A1 (nx65416), .A2 (nx66118)) ;
    and03 ix1533 (.Y (nx1532), .A0 (nx66160), .A1 (nx65416), .A2 (nx66058)) ;
    and03 ix1517 (.Y (nx1516), .A0 (nx66160), .A1 (nx65416), .A2 (nx66062)) ;
    and03 ix1483 (.Y (nx1482), .A0 (nx66160), .A1 (nx65416), .A2 (nx66066)) ;
    and03 ix1499 (.Y (nx1498), .A0 (nx66160), .A1 (nx65416), .A2 (nx66070)) ;
    and03 ix1463 (.Y (nx1462), .A0 (nx66160), .A1 (nx65416), .A2 (nx66074)) ;
    and03 ix1447 (.Y (nx1446), .A0 (nx66160), .A1 (nx65416), .A2 (nx66078)) ;
    and03 ix1413 (.Y (nx1412), .A0 (nx66162), .A1 (nx65418), .A2 (nx66082)) ;
    and03 ix1429 (.Y (nx1428), .A0 (nx66162), .A1 (nx65418), .A2 (nx66086)) ;
    and03 ix1391 (.Y (nx1390), .A0 (nx66162), .A1 (nx65418), .A2 (nx66090)) ;
    and03 ix1375 (.Y (nx1374), .A0 (nx66162), .A1 (nx65418), .A2 (nx66094)) ;
    and03 ix1341 (.Y (nx1340), .A0 (nx66162), .A1 (nx65418), .A2 (nx66098)) ;
    and03 ix1357 (.Y (nx1356), .A0 (nx66162), .A1 (nx65418), .A2 (nx66102)) ;
    and03 ix1321 (.Y (nx1320), .A0 (nx66162), .A1 (nx65418), .A2 (nx66106)) ;
    and03 ix1305 (.Y (nx1304), .A0 (nx65212), .A1 (nx65420), .A2 (nx66110)) ;
    and03 ix1271 (.Y (nx1270), .A0 (nx65212), .A1 (nx65420), .A2 (nx66114)) ;
    and03 ix1287 (.Y (nx1286), .A0 (nx65212), .A1 (nx65420), .A2 (nx66118)) ;
    and03 ix1233 (.Y (nx1232), .A0 (nx66164), .A1 (nx65420), .A2 (nx64524)) ;
    nor02ii ix55274 (.Y (nx55273), .A0 (address[6]), .A1 (address[7])) ;
    and03 ix1217 (.Y (nx1216), .A0 (nx66164), .A1 (nx65420), .A2 (nx64562)) ;
    and03 ix1183 (.Y (nx1182), .A0 (nx66164), .A1 (nx65420), .A2 (nx64600)) ;
    and03 ix1199 (.Y (nx1198), .A0 (nx66164), .A1 (nx65420), .A2 (nx64638)) ;
    and03 ix1163 (.Y (nx1162), .A0 (nx66164), .A1 (nx65422), .A2 (nx64676)) ;
    and03 ix1147 (.Y (nx1146), .A0 (nx66164), .A1 (nx65422), .A2 (nx64714)) ;
    and03 ix1113 (.Y (nx1112), .A0 (nx66166), .A1 (nx65422), .A2 (nx64752)) ;
    and03 ix1129 (.Y (nx1128), .A0 (nx66166), .A1 (nx65422), .A2 (nx64790)) ;
    and03 ix1091 (.Y (nx1090), .A0 (nx66166), .A1 (nx65422), .A2 (nx64828)) ;
    and03 ix1075 (.Y (nx1074), .A0 (nx66166), .A1 (nx65422), .A2 (nx64866)) ;
    and03 ix1041 (.Y (nx1040), .A0 (nx66166), .A1 (nx65422), .A2 (nx64904)) ;
    and03 ix1057 (.Y (nx1056), .A0 (nx66166), .A1 (nx65424), .A2 (nx64942)) ;
    and03 ix1021 (.Y (nx1020), .A0 (nx66166), .A1 (nx65424), .A2 (nx64980)) ;
    and03 ix1005 (.Y (nx1004), .A0 (nx65216), .A1 (nx65424), .A2 (nx65018)) ;
    and03 ix971 (.Y (nx970), .A0 (nx65216), .A1 (nx65424), .A2 (nx65056)) ;
    and03 ix987 (.Y (nx986), .A0 (nx65216), .A1 (nx65424), .A2 (nx65094)) ;
    and03 ix939 (.Y (nx938), .A0 (nx66168), .A1 (nx65424), .A2 (nx64524)) ;
    and03 ix923 (.Y (nx922), .A0 (nx66168), .A1 (nx65424), .A2 (nx64562)) ;
    and03 ix889 (.Y (nx888), .A0 (nx66168), .A1 (nx65426), .A2 (nx64600)) ;
    and03 ix905 (.Y (nx904), .A0 (nx66168), .A1 (nx65426), .A2 (nx64638)) ;
    and03 ix869 (.Y (nx868), .A0 (nx66168), .A1 (nx65426), .A2 (nx64676)) ;
    and03 ix853 (.Y (nx852), .A0 (nx66168), .A1 (nx65426), .A2 (nx64714)) ;
    and03 ix819 (.Y (nx818), .A0 (nx66170), .A1 (nx65426), .A2 (nx64752)) ;
    and03 ix835 (.Y (nx834), .A0 (nx66170), .A1 (nx65426), .A2 (nx64790)) ;
    and03 ix797 (.Y (nx796), .A0 (nx66170), .A1 (nx65426), .A2 (nx64828)) ;
    and03 ix781 (.Y (nx780), .A0 (nx66170), .A1 (nx65428), .A2 (nx64866)) ;
    and03 ix747 (.Y (nx746), .A0 (nx66170), .A1 (nx65428), .A2 (nx64904)) ;
    and03 ix763 (.Y (nx762), .A0 (nx66170), .A1 (nx65428), .A2 (nx64942)) ;
    and03 ix727 (.Y (nx726), .A0 (nx66170), .A1 (nx65428), .A2 (nx64980)) ;
    and03 ix711 (.Y (nx710), .A0 (nx65220), .A1 (nx65428), .A2 (nx65018)) ;
    and03 ix677 (.Y (nx676), .A0 (nx65220), .A1 (nx65428), .A2 (nx65056)) ;
    and03 ix693 (.Y (nx692), .A0 (nx65220), .A1 (nx65428), .A2 (nx65094)) ;
    and03 ix641 (.Y (nx640), .A0 (nx66172), .A1 (nx65430), .A2 (nx64524)) ;
    and03 ix625 (.Y (nx624), .A0 (nx66172), .A1 (nx65430), .A2 (nx64562)) ;
    and03 ix591 (.Y (nx590), .A0 (nx66172), .A1 (nx65430), .A2 (nx64600)) ;
    and03 ix607 (.Y (nx606), .A0 (nx66172), .A1 (nx65430), .A2 (nx64638)) ;
    and03 ix571 (.Y (nx570), .A0 (nx66172), .A1 (nx65430), .A2 (nx64676)) ;
    and03 ix555 (.Y (nx554), .A0 (nx66172), .A1 (nx65430), .A2 (nx64714)) ;
    and03 ix521 (.Y (nx520), .A0 (nx66174), .A1 (nx65430), .A2 (nx64752)) ;
    and03 ix537 (.Y (nx536), .A0 (nx66174), .A1 (nx65432), .A2 (nx64790)) ;
    and03 ix499 (.Y (nx498), .A0 (nx66174), .A1 (nx65432), .A2 (nx64828)) ;
    and03 ix483 (.Y (nx482), .A0 (nx66174), .A1 (nx65432), .A2 (nx64866)) ;
    and03 ix449 (.Y (nx448), .A0 (nx66174), .A1 (nx65432), .A2 (nx64904)) ;
    and03 ix465 (.Y (nx464), .A0 (nx66174), .A1 (nx65432), .A2 (nx64942)) ;
    and03 ix429 (.Y (nx428), .A0 (nx66174), .A1 (nx65432), .A2 (nx64980)) ;
    and03 ix413 (.Y (nx412), .A0 (nx65224), .A1 (nx65432), .A2 (nx65018)) ;
    and03 ix379 (.Y (nx378), .A0 (nx65224), .A1 (nx65434), .A2 (nx65056)) ;
    and03 ix395 (.Y (nx394), .A0 (nx65224), .A1 (nx65434), .A2 (nx65094)) ;
    and03 ix345 (.Y (nx344), .A0 (nx66176), .A1 (nx65434), .A2 (nx64524)) ;
    and03 ix327 (.Y (nx326), .A0 (nx66176), .A1 (nx65434), .A2 (nx64562)) ;
    and03 ix289 (.Y (nx288), .A0 (nx66176), .A1 (nx65434), .A2 (nx64600)) ;
    and03 ix307 (.Y (nx306), .A0 (nx66176), .A1 (nx65434), .A2 (nx64638)) ;
    and03 ix265 (.Y (nx264), .A0 (nx66176), .A1 (nx65434), .A2 (nx64676)) ;
    and03 ix247 (.Y (nx246), .A0 (nx66176), .A1 (nx65436), .A2 (nx64714)) ;
    and03 ix209 (.Y (nx208), .A0 (nx66178), .A1 (nx65436), .A2 (nx64752)) ;
    and03 ix227 (.Y (nx226), .A0 (nx66178), .A1 (nx65436), .A2 (nx64790)) ;
    and03 ix181 (.Y (nx180), .A0 (nx66178), .A1 (nx65436), .A2 (nx64828)) ;
    and03 ix163 (.Y (nx162), .A0 (nx66178), .A1 (nx65436), .A2 (nx64866)) ;
    and03 ix125 (.Y (nx124), .A0 (nx66178), .A1 (nx65436), .A2 (nx64904)) ;
    and03 ix143 (.Y (nx142), .A0 (nx66178), .A1 (nx65436), .A2 (nx64942)) ;
    and03 ix99 (.Y (nx98), .A0 (nx66178), .A1 (nx65438), .A2 (nx64980)) ;
    and03 ix79 (.Y (nx78), .A0 (nx65228), .A1 (nx65438), .A2 (nx65018)) ;
    and03 ix33 (.Y (nx32), .A0 (nx65228), .A1 (nx65438), .A2 (nx65056)) ;
    and03 ix55 (.Y (nx54), .A0 (nx65228), .A1 (nx65438), .A2 (nx65094)) ;
    inv02 ix65365 (.Y (nx65366), .A (nx66180)) ;
    inv02 ix65367 (.Y (nx65368), .A (nx66180)) ;
    inv02 ix65369 (.Y (nx65370), .A (nx66180)) ;
    inv02 ix65371 (.Y (nx65372), .A (nx66180)) ;
    inv02 ix65373 (.Y (nx65374), .A (nx66180)) ;
    inv02 ix65375 (.Y (nx65376), .A (nx66180)) ;
    inv02 ix65377 (.Y (nx65378), .A (nx66180)) ;
    inv02 ix65379 (.Y (nx65380), .A (nx66182)) ;
    inv02 ix65381 (.Y (nx65382), .A (nx66182)) ;
    inv02 ix65383 (.Y (nx65384), .A (nx66182)) ;
    inv02 ix65385 (.Y (nx65386), .A (nx66182)) ;
    inv02 ix65387 (.Y (nx65388), .A (nx66182)) ;
    inv02 ix65389 (.Y (nx65390), .A (nx66182)) ;
    inv02 ix65391 (.Y (nx65392), .A (nx66182)) ;
    inv02 ix65393 (.Y (nx65394), .A (nx66184)) ;
    inv02 ix65395 (.Y (nx65396), .A (nx66184)) ;
    inv02 ix65397 (.Y (nx65398), .A (nx66184)) ;
    inv02 ix65399 (.Y (nx65400), .A (nx66184)) ;
    inv02 ix65401 (.Y (nx65402), .A (nx66184)) ;
    inv02 ix65403 (.Y (nx65404), .A (nx66184)) ;
    inv02 ix65405 (.Y (nx65406), .A (nx66184)) ;
    inv02 ix65407 (.Y (nx65408), .A (nx66186)) ;
    inv02 ix65409 (.Y (nx65410), .A (nx66186)) ;
    inv02 ix65411 (.Y (nx65412), .A (nx66186)) ;
    inv02 ix65413 (.Y (nx65414), .A (nx66186)) ;
    inv02 ix65415 (.Y (nx65416), .A (nx66186)) ;
    inv02 ix65417 (.Y (nx65418), .A (nx66186)) ;
    inv02 ix65419 (.Y (nx65420), .A (nx66186)) ;
    inv02 ix65421 (.Y (nx65422), .A (nx66188)) ;
    inv02 ix65423 (.Y (nx65424), .A (nx66188)) ;
    inv02 ix65425 (.Y (nx65426), .A (nx66188)) ;
    inv02 ix65427 (.Y (nx65428), .A (nx66188)) ;
    inv02 ix65429 (.Y (nx65430), .A (nx66188)) ;
    inv02 ix65431 (.Y (nx65432), .A (nx66188)) ;
    inv02 ix65433 (.Y (nx65434), .A (nx66188)) ;
    inv02 ix65435 (.Y (nx65436), .A (nx66190)) ;
    inv02 ix65437 (.Y (nx65438), .A (nx66190)) ;
    buf02 ix65439 (.Y (nx65440), .A (address[5])) ;
    buf02 ix65441 (.Y (nx65442), .A (address[5])) ;
    buf02 ix65443 (.Y (nx65444), .A (address[1])) ;
    buf02 ix65445 (.Y (nx65446), .A (address[1])) ;
    inv02 ix65449 (.Y (nx65450), .A (nx66192)) ;
    inv02 ix65451 (.Y (nx65452), .A (nx66192)) ;
    inv02 ix65453 (.Y (nx65454), .A (nx66192)) ;
    inv02 ix65455 (.Y (nx65456), .A (nx66192)) ;
    inv02 ix65457 (.Y (nx65458), .A (nx66192)) ;
    inv02 ix65459 (.Y (nx65460), .A (nx66192)) ;
    inv02 ix65461 (.Y (nx65462), .A (nx66192)) ;
    inv02 ix65463 (.Y (nx65464), .A (nx66194)) ;
    inv02 ix65465 (.Y (nx65466), .A (nx66194)) ;
    inv02 ix65467 (.Y (nx65468), .A (nx66194)) ;
    inv02 ix65469 (.Y (nx65470), .A (nx66194)) ;
    inv02 ix65471 (.Y (nx65472), .A (nx66194)) ;
    inv02 ix65473 (.Y (nx65474), .A (nx66194)) ;
    inv02 ix65475 (.Y (nx65476), .A (nx66194)) ;
    inv02 ix65477 (.Y (nx65478), .A (nx66196)) ;
    inv02 ix65479 (.Y (nx65480), .A (nx66196)) ;
    inv02 ix65481 (.Y (nx65482), .A (nx66196)) ;
    inv02 ix65483 (.Y (nx65484), .A (nx66196)) ;
    inv02 ix65485 (.Y (nx65486), .A (nx66196)) ;
    inv02 ix65487 (.Y (nx65488), .A (nx66196)) ;
    inv02 ix65489 (.Y (nx65490), .A (nx66196)) ;
    inv02 ix65491 (.Y (nx65492), .A (nx66198)) ;
    inv02 ix65493 (.Y (nx65494), .A (nx66198)) ;
    inv02 ix65495 (.Y (nx65496), .A (nx66198)) ;
    inv02 ix65497 (.Y (nx65498), .A (nx66198)) ;
    inv02 ix65499 (.Y (nx65500), .A (nx66198)) ;
    inv02 ix65501 (.Y (nx65502), .A (nx66198)) ;
    inv02 ix65503 (.Y (nx65504), .A (nx66198)) ;
    inv02 ix65505 (.Y (nx65506), .A (nx66200)) ;
    inv02 ix65507 (.Y (nx65508), .A (nx66200)) ;
    inv02 ix65509 (.Y (nx65510), .A (nx66200)) ;
    inv02 ix65511 (.Y (nx65512), .A (nx66200)) ;
    inv02 ix65513 (.Y (nx65514), .A (nx66200)) ;
    inv02 ix65515 (.Y (nx65516), .A (nx66200)) ;
    inv02 ix65517 (.Y (nx65518), .A (nx66200)) ;
    inv02 ix65519 (.Y (nx65520), .A (nx66202)) ;
    inv02 ix65521 (.Y (nx65522), .A (nx66202)) ;
    inv02 ix65525 (.Y (nx65526), .A (nx66204)) ;
    inv02 ix65527 (.Y (nx65528), .A (nx66204)) ;
    inv02 ix65529 (.Y (nx65530), .A (nx66204)) ;
    inv02 ix65531 (.Y (nx65532), .A (nx66204)) ;
    inv02 ix65533 (.Y (nx65534), .A (nx66204)) ;
    inv02 ix65535 (.Y (nx65536), .A (nx66204)) ;
    inv02 ix65537 (.Y (nx65538), .A (nx66204)) ;
    inv02 ix65539 (.Y (nx65540), .A (nx66206)) ;
    inv02 ix65541 (.Y (nx65542), .A (nx66206)) ;
    inv02 ix65543 (.Y (nx65544), .A (nx66206)) ;
    inv02 ix65545 (.Y (nx65546), .A (nx66206)) ;
    inv02 ix65547 (.Y (nx65548), .A (nx66206)) ;
    inv02 ix65549 (.Y (nx65550), .A (nx66206)) ;
    inv02 ix65551 (.Y (nx65552), .A (nx66206)) ;
    inv02 ix65553 (.Y (nx65554), .A (nx66208)) ;
    inv02 ix65555 (.Y (nx65556), .A (nx66208)) ;
    inv02 ix65557 (.Y (nx65558), .A (nx66208)) ;
    inv02 ix65559 (.Y (nx65560), .A (nx66208)) ;
    inv02 ix65561 (.Y (nx65562), .A (nx66208)) ;
    inv02 ix65563 (.Y (nx65564), .A (nx66208)) ;
    inv02 ix65565 (.Y (nx65566), .A (nx66208)) ;
    inv02 ix65567 (.Y (nx65568), .A (nx66210)) ;
    inv02 ix65569 (.Y (nx65570), .A (nx66210)) ;
    inv02 ix65571 (.Y (nx65572), .A (nx66210)) ;
    inv02 ix65573 (.Y (nx65574), .A (nx66210)) ;
    inv02 ix65575 (.Y (nx65576), .A (nx66210)) ;
    inv02 ix65577 (.Y (nx65578), .A (nx66210)) ;
    inv02 ix65579 (.Y (nx65580), .A (nx66210)) ;
    inv02 ix65581 (.Y (nx65582), .A (nx66212)) ;
    inv02 ix65583 (.Y (nx65584), .A (nx66212)) ;
    inv02 ix65585 (.Y (nx65586), .A (nx66212)) ;
    inv02 ix65587 (.Y (nx65588), .A (nx66212)) ;
    inv02 ix65589 (.Y (nx65590), .A (nx66212)) ;
    inv02 ix65591 (.Y (nx65592), .A (nx66212)) ;
    inv02 ix65593 (.Y (nx65594), .A (nx66212)) ;
    inv02 ix65595 (.Y (nx65596), .A (nx66214)) ;
    inv02 ix65597 (.Y (nx65598), .A (nx66214)) ;
    inv02 ix65601 (.Y (nx65602), .A (nx66216)) ;
    inv02 ix65603 (.Y (nx65604), .A (nx66216)) ;
    inv02 ix65605 (.Y (nx65606), .A (nx66216)) ;
    inv02 ix65607 (.Y (nx65608), .A (nx66216)) ;
    inv02 ix65609 (.Y (nx65610), .A (nx66216)) ;
    inv02 ix65611 (.Y (nx65612), .A (nx66216)) ;
    inv02 ix65613 (.Y (nx65614), .A (nx66216)) ;
    inv02 ix65615 (.Y (nx65616), .A (nx66218)) ;
    inv02 ix65617 (.Y (nx65618), .A (nx66218)) ;
    inv02 ix65619 (.Y (nx65620), .A (nx66218)) ;
    inv02 ix65621 (.Y (nx65622), .A (nx66218)) ;
    inv02 ix65623 (.Y (nx65624), .A (nx66218)) ;
    inv02 ix65625 (.Y (nx65626), .A (nx66218)) ;
    inv02 ix65627 (.Y (nx65628), .A (nx66218)) ;
    inv02 ix65629 (.Y (nx65630), .A (nx66220)) ;
    inv02 ix65631 (.Y (nx65632), .A (nx66220)) ;
    inv02 ix65633 (.Y (nx65634), .A (nx66220)) ;
    inv02 ix65635 (.Y (nx65636), .A (nx66220)) ;
    inv02 ix65637 (.Y (nx65638), .A (nx66220)) ;
    inv02 ix65639 (.Y (nx65640), .A (nx66220)) ;
    inv02 ix65641 (.Y (nx65642), .A (nx66220)) ;
    inv02 ix65643 (.Y (nx65644), .A (nx66222)) ;
    inv02 ix65645 (.Y (nx65646), .A (nx66222)) ;
    inv02 ix65647 (.Y (nx65648), .A (nx66222)) ;
    inv02 ix65649 (.Y (nx65650), .A (nx66222)) ;
    inv02 ix65651 (.Y (nx65652), .A (nx66222)) ;
    inv02 ix65653 (.Y (nx65654), .A (nx66222)) ;
    inv02 ix65655 (.Y (nx65656), .A (nx66222)) ;
    inv02 ix65657 (.Y (nx65658), .A (nx66224)) ;
    inv02 ix65659 (.Y (nx65660), .A (nx66224)) ;
    inv02 ix65661 (.Y (nx65662), .A (nx66224)) ;
    inv02 ix65663 (.Y (nx65664), .A (nx66224)) ;
    inv02 ix65665 (.Y (nx65666), .A (nx66224)) ;
    inv02 ix65667 (.Y (nx65668), .A (nx66224)) ;
    inv02 ix65669 (.Y (nx65670), .A (nx66224)) ;
    inv02 ix65671 (.Y (nx65672), .A (nx66226)) ;
    inv02 ix65673 (.Y (nx65674), .A (nx66226)) ;
    inv02 ix65677 (.Y (nx65678), .A (nx66228)) ;
    inv02 ix65679 (.Y (nx65680), .A (nx66228)) ;
    inv02 ix65681 (.Y (nx65682), .A (nx66228)) ;
    inv02 ix65683 (.Y (nx65684), .A (nx66228)) ;
    inv02 ix65685 (.Y (nx65686), .A (nx66228)) ;
    inv02 ix65687 (.Y (nx65688), .A (nx66228)) ;
    inv02 ix65689 (.Y (nx65690), .A (nx66228)) ;
    inv02 ix65691 (.Y (nx65692), .A (nx66230)) ;
    inv02 ix65693 (.Y (nx65694), .A (nx66230)) ;
    inv02 ix65695 (.Y (nx65696), .A (nx66230)) ;
    inv02 ix65697 (.Y (nx65698), .A (nx66230)) ;
    inv02 ix65699 (.Y (nx65700), .A (nx66230)) ;
    inv02 ix65701 (.Y (nx65702), .A (nx66230)) ;
    inv02 ix65703 (.Y (nx65704), .A (nx66230)) ;
    inv02 ix65705 (.Y (nx65706), .A (nx66232)) ;
    inv02 ix65707 (.Y (nx65708), .A (nx66232)) ;
    inv02 ix65709 (.Y (nx65710), .A (nx66232)) ;
    inv02 ix65711 (.Y (nx65712), .A (nx66232)) ;
    inv02 ix65713 (.Y (nx65714), .A (nx66232)) ;
    inv02 ix65715 (.Y (nx65716), .A (nx66232)) ;
    inv02 ix65717 (.Y (nx65718), .A (nx66232)) ;
    inv02 ix65719 (.Y (nx65720), .A (nx66234)) ;
    inv02 ix65721 (.Y (nx65722), .A (nx66234)) ;
    inv02 ix65723 (.Y (nx65724), .A (nx66234)) ;
    inv02 ix65725 (.Y (nx65726), .A (nx66234)) ;
    inv02 ix65727 (.Y (nx65728), .A (nx66234)) ;
    inv02 ix65729 (.Y (nx65730), .A (nx66234)) ;
    inv02 ix65731 (.Y (nx65732), .A (nx66234)) ;
    inv02 ix65733 (.Y (nx65734), .A (nx66236)) ;
    inv02 ix65735 (.Y (nx65736), .A (nx66236)) ;
    inv02 ix65737 (.Y (nx65738), .A (nx66236)) ;
    inv02 ix65739 (.Y (nx65740), .A (nx66236)) ;
    inv02 ix65741 (.Y (nx65742), .A (nx66236)) ;
    inv02 ix65743 (.Y (nx65744), .A (nx66236)) ;
    inv02 ix65745 (.Y (nx65746), .A (nx66236)) ;
    inv02 ix65747 (.Y (nx65748), .A (nx66238)) ;
    inv02 ix65749 (.Y (nx65750), .A (nx66238)) ;
    inv02 ix65753 (.Y (nx65754), .A (nx66240)) ;
    inv02 ix65755 (.Y (nx65756), .A (nx66240)) ;
    inv02 ix65757 (.Y (nx65758), .A (nx66240)) ;
    inv02 ix65759 (.Y (nx65760), .A (nx66240)) ;
    inv02 ix65761 (.Y (nx65762), .A (nx66240)) ;
    inv02 ix65763 (.Y (nx65764), .A (nx66240)) ;
    inv02 ix65765 (.Y (nx65766), .A (nx66240)) ;
    inv02 ix65767 (.Y (nx65768), .A (nx66242)) ;
    inv02 ix65769 (.Y (nx65770), .A (nx66242)) ;
    inv02 ix65771 (.Y (nx65772), .A (nx66242)) ;
    inv02 ix65773 (.Y (nx65774), .A (nx66242)) ;
    inv02 ix65775 (.Y (nx65776), .A (nx66242)) ;
    inv02 ix65777 (.Y (nx65778), .A (nx66242)) ;
    inv02 ix65779 (.Y (nx65780), .A (nx66242)) ;
    inv02 ix65781 (.Y (nx65782), .A (nx66244)) ;
    inv02 ix65783 (.Y (nx65784), .A (nx66244)) ;
    inv02 ix65785 (.Y (nx65786), .A (nx66244)) ;
    inv02 ix65787 (.Y (nx65788), .A (nx66244)) ;
    inv02 ix65789 (.Y (nx65790), .A (nx66244)) ;
    inv02 ix65791 (.Y (nx65792), .A (nx66244)) ;
    inv02 ix65793 (.Y (nx65794), .A (nx66244)) ;
    inv02 ix65795 (.Y (nx65796), .A (nx66246)) ;
    inv02 ix65797 (.Y (nx65798), .A (nx66246)) ;
    inv02 ix65799 (.Y (nx65800), .A (nx66246)) ;
    inv02 ix65801 (.Y (nx65802), .A (nx66246)) ;
    inv02 ix65803 (.Y (nx65804), .A (nx66246)) ;
    inv02 ix65805 (.Y (nx65806), .A (nx66246)) ;
    inv02 ix65807 (.Y (nx65808), .A (nx66246)) ;
    inv02 ix65809 (.Y (nx65810), .A (nx66248)) ;
    inv02 ix65811 (.Y (nx65812), .A (nx66248)) ;
    inv02 ix65813 (.Y (nx65814), .A (nx66248)) ;
    inv02 ix65815 (.Y (nx65816), .A (nx66248)) ;
    inv02 ix65817 (.Y (nx65818), .A (nx66248)) ;
    inv02 ix65819 (.Y (nx65820), .A (nx66248)) ;
    inv02 ix65821 (.Y (nx65822), .A (nx66248)) ;
    inv02 ix65823 (.Y (nx65824), .A (nx66250)) ;
    inv02 ix65825 (.Y (nx65826), .A (nx66250)) ;
    inv02 ix65829 (.Y (nx65830), .A (nx66252)) ;
    inv02 ix65831 (.Y (nx65832), .A (nx66252)) ;
    inv02 ix65833 (.Y (nx65834), .A (nx66252)) ;
    inv02 ix65835 (.Y (nx65836), .A (nx66252)) ;
    inv02 ix65837 (.Y (nx65838), .A (nx66252)) ;
    inv02 ix65839 (.Y (nx65840), .A (nx66252)) ;
    inv02 ix65841 (.Y (nx65842), .A (nx66252)) ;
    inv02 ix65843 (.Y (nx65844), .A (nx66254)) ;
    inv02 ix65845 (.Y (nx65846), .A (nx66254)) ;
    inv02 ix65847 (.Y (nx65848), .A (nx66254)) ;
    inv02 ix65849 (.Y (nx65850), .A (nx66254)) ;
    inv02 ix65851 (.Y (nx65852), .A (nx66254)) ;
    inv02 ix65853 (.Y (nx65854), .A (nx66254)) ;
    inv02 ix65855 (.Y (nx65856), .A (nx66254)) ;
    inv02 ix65857 (.Y (nx65858), .A (nx66256)) ;
    inv02 ix65859 (.Y (nx65860), .A (nx66256)) ;
    inv02 ix65861 (.Y (nx65862), .A (nx66256)) ;
    inv02 ix65863 (.Y (nx65864), .A (nx66256)) ;
    inv02 ix65865 (.Y (nx65866), .A (nx66256)) ;
    inv02 ix65867 (.Y (nx65868), .A (nx66256)) ;
    inv02 ix65869 (.Y (nx65870), .A (nx66256)) ;
    inv02 ix65871 (.Y (nx65872), .A (nx66258)) ;
    inv02 ix65873 (.Y (nx65874), .A (nx66258)) ;
    inv02 ix65875 (.Y (nx65876), .A (nx66258)) ;
    inv02 ix65877 (.Y (nx65878), .A (nx66258)) ;
    inv02 ix65879 (.Y (nx65880), .A (nx66258)) ;
    inv02 ix65881 (.Y (nx65882), .A (nx66258)) ;
    inv02 ix65883 (.Y (nx65884), .A (nx66258)) ;
    inv02 ix65885 (.Y (nx65886), .A (nx66260)) ;
    inv02 ix65887 (.Y (nx65888), .A (nx66260)) ;
    inv02 ix65889 (.Y (nx65890), .A (nx66260)) ;
    inv02 ix65891 (.Y (nx65892), .A (nx66260)) ;
    inv02 ix65893 (.Y (nx65894), .A (nx66260)) ;
    inv02 ix65895 (.Y (nx65896), .A (nx66260)) ;
    inv02 ix65897 (.Y (nx65898), .A (nx66260)) ;
    inv02 ix65899 (.Y (nx65900), .A (nx66262)) ;
    inv02 ix65901 (.Y (nx65902), .A (nx66262)) ;
    inv02 ix65905 (.Y (nx65906), .A (nx66264)) ;
    inv02 ix65907 (.Y (nx65908), .A (nx66264)) ;
    inv02 ix65909 (.Y (nx65910), .A (nx66264)) ;
    inv02 ix65911 (.Y (nx65912), .A (nx66264)) ;
    inv02 ix65913 (.Y (nx65914), .A (nx66264)) ;
    inv02 ix65915 (.Y (nx65916), .A (nx66264)) ;
    inv02 ix65917 (.Y (nx65918), .A (nx66264)) ;
    inv02 ix65919 (.Y (nx65920), .A (nx66266)) ;
    inv02 ix65921 (.Y (nx65922), .A (nx66266)) ;
    inv02 ix65923 (.Y (nx65924), .A (nx66266)) ;
    inv02 ix65925 (.Y (nx65926), .A (nx66266)) ;
    inv02 ix65927 (.Y (nx65928), .A (nx66266)) ;
    inv02 ix65929 (.Y (nx65930), .A (nx66266)) ;
    inv02 ix65931 (.Y (nx65932), .A (nx66266)) ;
    inv02 ix65933 (.Y (nx65934), .A (nx66268)) ;
    inv02 ix65935 (.Y (nx65936), .A (nx66268)) ;
    inv02 ix65937 (.Y (nx65938), .A (nx66268)) ;
    inv02 ix65939 (.Y (nx65940), .A (nx66268)) ;
    inv02 ix65941 (.Y (nx65942), .A (nx66268)) ;
    inv02 ix65943 (.Y (nx65944), .A (nx66268)) ;
    inv02 ix65945 (.Y (nx65946), .A (nx66268)) ;
    inv02 ix65947 (.Y (nx65948), .A (nx66270)) ;
    inv02 ix65949 (.Y (nx65950), .A (nx66270)) ;
    inv02 ix65951 (.Y (nx65952), .A (nx66270)) ;
    inv02 ix65953 (.Y (nx65954), .A (nx66270)) ;
    inv02 ix65955 (.Y (nx65956), .A (nx66270)) ;
    inv02 ix65957 (.Y (nx65958), .A (nx66270)) ;
    inv02 ix65959 (.Y (nx65960), .A (nx66270)) ;
    inv02 ix65961 (.Y (nx65962), .A (nx66272)) ;
    inv02 ix65963 (.Y (nx65964), .A (nx66272)) ;
    inv02 ix65965 (.Y (nx65966), .A (nx66272)) ;
    inv02 ix65967 (.Y (nx65968), .A (nx66272)) ;
    inv02 ix65969 (.Y (nx65970), .A (nx66272)) ;
    inv02 ix65971 (.Y (nx65972), .A (nx66272)) ;
    inv02 ix65973 (.Y (nx65974), .A (nx66272)) ;
    inv02 ix65975 (.Y (nx65976), .A (nx66274)) ;
    inv02 ix65977 (.Y (nx65978), .A (nx66274)) ;
    inv02 ix65981 (.Y (nx65982), .A (nx66276)) ;
    inv02 ix65983 (.Y (nx65984), .A (nx66276)) ;
    inv02 ix65985 (.Y (nx65986), .A (nx66276)) ;
    inv02 ix65987 (.Y (nx65988), .A (nx66276)) ;
    inv02 ix65989 (.Y (nx65990), .A (nx66276)) ;
    inv02 ix65991 (.Y (nx65992), .A (nx66276)) ;
    inv02 ix65993 (.Y (nx65994), .A (nx66276)) ;
    inv02 ix65995 (.Y (nx65996), .A (nx66278)) ;
    inv02 ix65997 (.Y (nx65998), .A (nx66278)) ;
    inv02 ix65999 (.Y (nx66000), .A (nx66278)) ;
    inv02 ix66001 (.Y (nx66002), .A (nx66278)) ;
    inv02 ix66003 (.Y (nx66004), .A (nx66278)) ;
    inv02 ix66005 (.Y (nx66006), .A (nx66278)) ;
    inv02 ix66007 (.Y (nx66008), .A (nx66278)) ;
    inv02 ix66009 (.Y (nx66010), .A (nx66280)) ;
    inv02 ix66011 (.Y (nx66012), .A (nx66280)) ;
    inv02 ix66013 (.Y (nx66014), .A (nx66280)) ;
    inv02 ix66015 (.Y (nx66016), .A (nx66280)) ;
    inv02 ix66017 (.Y (nx66018), .A (nx66280)) ;
    inv02 ix66019 (.Y (nx66020), .A (nx66280)) ;
    inv02 ix66021 (.Y (nx66022), .A (nx66280)) ;
    inv02 ix66023 (.Y (nx66024), .A (nx66282)) ;
    inv02 ix66025 (.Y (nx66026), .A (nx66282)) ;
    inv02 ix66027 (.Y (nx66028), .A (nx66282)) ;
    inv02 ix66029 (.Y (nx66030), .A (nx66282)) ;
    inv02 ix66031 (.Y (nx66032), .A (nx66282)) ;
    inv02 ix66033 (.Y (nx66034), .A (nx66282)) ;
    inv02 ix66035 (.Y (nx66036), .A (nx66282)) ;
    inv02 ix66037 (.Y (nx66038), .A (nx66284)) ;
    inv02 ix66039 (.Y (nx66040), .A (nx66284)) ;
    inv02 ix66041 (.Y (nx66042), .A (nx66284)) ;
    inv02 ix66043 (.Y (nx66044), .A (nx66284)) ;
    inv02 ix66045 (.Y (nx66046), .A (nx66284)) ;
    inv02 ix66047 (.Y (nx66048), .A (nx66284)) ;
    inv02 ix66049 (.Y (nx66050), .A (nx66284)) ;
    inv02 ix66051 (.Y (nx66052), .A (nx66286)) ;
    inv02 ix66053 (.Y (nx66054), .A (nx66286)) ;
    inv02 ix66055 (.Y (nx66056), .A (nx65328)) ;
    inv02 ix66057 (.Y (nx66058), .A (nx65328)) ;
    inv02 ix66059 (.Y (nx66060), .A (nx65322)) ;
    inv02 ix66061 (.Y (nx66062), .A (nx65322)) ;
    inv02 ix66063 (.Y (nx66064), .A (nx65310)) ;
    inv02 ix66065 (.Y (nx66066), .A (nx65310)) ;
    inv02 ix66067 (.Y (nx66068), .A (nx65316)) ;
    inv02 ix66069 (.Y (nx66070), .A (nx65316)) ;
    inv02 ix66071 (.Y (nx66072), .A (nx65304)) ;
    inv02 ix66073 (.Y (nx66074), .A (nx65304)) ;
    inv02 ix66075 (.Y (nx66076), .A (nx65298)) ;
    inv02 ix66077 (.Y (nx66078), .A (nx65298)) ;
    inv02 ix66079 (.Y (nx66080), .A (nx65286)) ;
    inv02 ix66081 (.Y (nx66082), .A (nx65286)) ;
    inv02 ix66083 (.Y (nx66084), .A (nx65292)) ;
    inv02 ix66085 (.Y (nx66086), .A (nx65292)) ;
    inv02 ix66087 (.Y (nx66088), .A (nx65280)) ;
    inv02 ix66089 (.Y (nx66090), .A (nx65280)) ;
    inv02 ix66091 (.Y (nx66092), .A (nx65274)) ;
    inv02 ix66093 (.Y (nx66094), .A (nx65274)) ;
    inv02 ix66095 (.Y (nx66096), .A (nx65262)) ;
    inv02 ix66097 (.Y (nx66098), .A (nx65262)) ;
    inv02 ix66099 (.Y (nx66100), .A (nx65268)) ;
    inv02 ix66101 (.Y (nx66102), .A (nx65268)) ;
    inv02 ix66103 (.Y (nx66104), .A (nx65256)) ;
    inv02 ix66105 (.Y (nx66106), .A (nx65256)) ;
    inv02 ix66107 (.Y (nx66108), .A (nx65250)) ;
    inv02 ix66109 (.Y (nx66110), .A (nx65250)) ;
    inv02 ix66111 (.Y (nx66112), .A (nx65238)) ;
    inv02 ix66113 (.Y (nx66114), .A (nx65238)) ;
    inv02 ix66115 (.Y (nx66116), .A (nx65244)) ;
    inv02 ix66117 (.Y (nx66118), .A (nx65244)) ;
    inv02 ix66119 (.Y (nx66120), .A (nx4498)) ;
    inv02 ix66121 (.Y (nx66122), .A (nx4498)) ;
    inv02 ix66123 (.Y (nx66124), .A (nx4206)) ;
    inv02 ix66125 (.Y (nx66126), .A (nx4206)) ;
    inv02 ix66127 (.Y (nx66128), .A (nx3912)) ;
    inv02 ix66129 (.Y (nx66130), .A (nx3912)) ;
    inv02 ix66131 (.Y (nx66132), .A (nx3620)) ;
    inv02 ix66133 (.Y (nx66134), .A (nx3620)) ;
    inv02 ix66135 (.Y (nx66136), .A (nx3318)) ;
    inv02 ix66137 (.Y (nx66138), .A (nx3318)) ;
    inv02 ix66139 (.Y (nx66140), .A (nx3026)) ;
    inv02 ix66141 (.Y (nx66142), .A (nx3026)) ;
    inv02 ix66143 (.Y (nx66144), .A (nx2732)) ;
    inv02 ix66145 (.Y (nx66146), .A (nx2732)) ;
    inv02 ix66147 (.Y (nx66148), .A (nx2440)) ;
    inv02 ix66149 (.Y (nx66150), .A (nx2440)) ;
    inv02 ix66151 (.Y (nx66152), .A (nx2142)) ;
    inv02 ix66153 (.Y (nx66154), .A (nx2142)) ;
    inv02 ix66155 (.Y (nx66156), .A (nx1554)) ;
    inv02 ix66157 (.Y (nx66158), .A (nx1554)) ;
    inv02 ix66159 (.Y (nx66160), .A (nx1262)) ;
    inv02 ix66161 (.Y (nx66162), .A (nx1262)) ;
    inv02 ix66163 (.Y (nx66164), .A (nx962)) ;
    inv02 ix66165 (.Y (nx66166), .A (nx962)) ;
    inv02 ix66167 (.Y (nx66168), .A (nx668)) ;
    inv02 ix66169 (.Y (nx66170), .A (nx668)) ;
    inv02 ix66171 (.Y (nx66172), .A (nx370)) ;
    inv02 ix66173 (.Y (nx66174), .A (nx370)) ;
    inv02 ix66175 (.Y (nx66176), .A (nx10)) ;
    inv02 ix66177 (.Y (nx66178), .A (nx10)) ;
    inv02 ix66179 (.Y (nx66180), .A (write_en)) ;
    inv02 ix66181 (.Y (nx66182), .A (write_en)) ;
    inv02 ix66183 (.Y (nx66184), .A (write_en)) ;
    inv02 ix66185 (.Y (nx66186), .A (write_en)) ;
    inv02 ix66187 (.Y (nx66188), .A (write_en)) ;
    inv02 ix66189 (.Y (nx66190), .A (write_en)) ;
    inv02 ix66191 (.Y (nx66192), .A (datain[7])) ;
    inv02 ix66193 (.Y (nx66194), .A (datain[7])) ;
    inv02 ix66195 (.Y (nx66196), .A (datain[7])) ;
    inv02 ix66197 (.Y (nx66198), .A (datain[7])) ;
    inv02 ix66199 (.Y (nx66200), .A (datain[7])) ;
    inv02 ix66201 (.Y (nx66202), .A (datain[7])) ;
    inv02 ix66203 (.Y (nx66204), .A (datain[6])) ;
    inv02 ix66205 (.Y (nx66206), .A (datain[6])) ;
    inv02 ix66207 (.Y (nx66208), .A (datain[6])) ;
    inv02 ix66209 (.Y (nx66210), .A (datain[6])) ;
    inv02 ix66211 (.Y (nx66212), .A (datain[6])) ;
    inv02 ix66213 (.Y (nx66214), .A (datain[6])) ;
    inv02 ix66215 (.Y (nx66216), .A (datain[5])) ;
    inv02 ix66217 (.Y (nx66218), .A (datain[5])) ;
    inv02 ix66219 (.Y (nx66220), .A (datain[5])) ;
    inv02 ix66221 (.Y (nx66222), .A (datain[5])) ;
    inv02 ix66223 (.Y (nx66224), .A (datain[5])) ;
    inv02 ix66225 (.Y (nx66226), .A (datain[5])) ;
    inv02 ix66227 (.Y (nx66228), .A (datain[4])) ;
    inv02 ix66229 (.Y (nx66230), .A (datain[4])) ;
    inv02 ix66231 (.Y (nx66232), .A (datain[4])) ;
    inv02 ix66233 (.Y (nx66234), .A (datain[4])) ;
    inv02 ix66235 (.Y (nx66236), .A (datain[4])) ;
    inv02 ix66237 (.Y (nx66238), .A (datain[4])) ;
    inv02 ix66239 (.Y (nx66240), .A (datain[3])) ;
    inv02 ix66241 (.Y (nx66242), .A (datain[3])) ;
    inv02 ix66243 (.Y (nx66244), .A (datain[3])) ;
    inv02 ix66245 (.Y (nx66246), .A (datain[3])) ;
    inv02 ix66247 (.Y (nx66248), .A (datain[3])) ;
    inv02 ix66249 (.Y (nx66250), .A (datain[3])) ;
    inv02 ix66251 (.Y (nx66252), .A (datain[2])) ;
    inv02 ix66253 (.Y (nx66254), .A (datain[2])) ;
    inv02 ix66255 (.Y (nx66256), .A (datain[2])) ;
    inv02 ix66257 (.Y (nx66258), .A (datain[2])) ;
    inv02 ix66259 (.Y (nx66260), .A (datain[2])) ;
    inv02 ix66261 (.Y (nx66262), .A (datain[2])) ;
    inv02 ix66263 (.Y (nx66264), .A (datain[1])) ;
    inv02 ix66265 (.Y (nx66266), .A (datain[1])) ;
    inv02 ix66267 (.Y (nx66268), .A (datain[1])) ;
    inv02 ix66269 (.Y (nx66270), .A (datain[1])) ;
    inv02 ix66271 (.Y (nx66272), .A (datain[1])) ;
    inv02 ix66273 (.Y (nx66274), .A (datain[1])) ;
    inv02 ix66275 (.Y (nx66276), .A (datain[0])) ;
    inv02 ix66277 (.Y (nx66278), .A (datain[0])) ;
    inv02 ix66279 (.Y (nx66280), .A (datain[0])) ;
    inv02 ix66281 (.Y (nx66282), .A (datain[0])) ;
    inv02 ix66283 (.Y (nx66284), .A (datain[0])) ;
    inv02 ix66285 (.Y (nx66286), .A (datain[0])) ;
endmodule


module nbit_mux2x1_8 ( input1, input2, s0, \output  ) ;

    input [7:0]input1 ;
    input [7:0]input2 ;
    input s0 ;
    output [7:0]\output  ;

    wire nx157, nx159;



    mux21_ni ix7 (.Y (\output [0]), .A0 (input1[0]), .A1 (input2[0]), .S0 (nx157
             )) ;
    mux21_ni ix15 (.Y (\output [1]), .A0 (input1[1]), .A1 (input2[1]), .S0 (
             nx157)) ;
    mux21_ni ix23 (.Y (\output [2]), .A0 (input1[2]), .A1 (input2[2]), .S0 (
             nx157)) ;
    mux21_ni ix31 (.Y (\output [3]), .A0 (input1[3]), .A1 (input2[3]), .S0 (
             nx157)) ;
    mux21_ni ix39 (.Y (\output [4]), .A0 (input1[4]), .A1 (input2[4]), .S0 (
             nx157)) ;
    mux21_ni ix47 (.Y (\output [5]), .A0 (input1[5]), .A1 (input2[5]), .S0 (
             nx157)) ;
    mux21_ni ix55 (.Y (\output [6]), .A0 (input1[6]), .A1 (input2[6]), .S0 (
             nx157)) ;
    mux21_ni ix63 (.Y (\output [7]), .A0 (input1[7]), .A1 (input2[7]), .S0 (
             nx159)) ;
    buf02 ix156 (.Y (nx157), .A (s0)) ;
    buf02 ix158 (.Y (nx159), .A (s0)) ;
endmodule

