//
// Verilog description for cell system, 
// Sat May 13 10:16:06 2017
//
// LeonardoSpectrum Level 3, 2016a.6 
//


module system ( clk, rst, start, motor_done, nvm_input_address, zero, one, done, 
                motor_move, motor_direction ) ;

    input clk ;
    input rst ;
    input start ;
    input motor_done ;
    input [11:0]nvm_input_address ;
    input zero ;
    input one ;
    output done ;
    output motor_move ;
    output [0:0]motor_direction ;

    wire nvm_data_127, nvm_data_126, nvm_data_125, nvm_data_124, nvm_data_123, 
         nvm_data_122, nvm_data_121, nvm_data_120, nvm_data_119, nvm_data_118, 
         nvm_data_117, nvm_data_116, nvm_data_115, nvm_data_114, nvm_data_113, 
         nvm_data_112, nvm_data_111, nvm_data_110, nvm_data_109, nvm_data_108, 
         nvm_data_107, nvm_data_106, nvm_data_105, nvm_data_104, nvm_data_103, 
         nvm_data_102, nvm_data_101, nvm_data_100, nvm_data_99, nvm_data_98, 
         nvm_data_97, nvm_data_96, nvm_data_95, nvm_data_94, nvm_data_93, 
         nvm_data_92, nvm_data_91, nvm_data_90, nvm_data_89, nvm_data_88, 
         nvm_data_87, nvm_data_86, nvm_data_85, nvm_data_84, nvm_data_83, 
         nvm_data_82, nvm_data_81, nvm_data_80, nvm_data_79, nvm_data_78, 
         nvm_data_77, nvm_data_76, nvm_data_75, nvm_data_74, nvm_data_73, 
         nvm_data_72, nvm_data_71, nvm_data_70, nvm_data_69, nvm_data_68, 
         nvm_data_67, nvm_data_66, nvm_data_65, nvm_data_64, nvm_data_63, 
         nvm_data_62, nvm_data_61, nvm_data_60, nvm_data_59, nvm_data_58, 
         nvm_data_57, nvm_data_56, nvm_data_55, nvm_data_54, nvm_data_53, 
         nvm_data_52, nvm_data_51, nvm_data_50, nvm_data_49, nvm_data_48, 
         nvm_data_47, nvm_data_46, nvm_data_45, nvm_data_44, nvm_data_43, 
         nvm_data_42, nvm_data_41, nvm_data_40, nvm_data_39, nvm_data_38, 
         nvm_data_37, nvm_data_36, nvm_data_35, nvm_data_34, nvm_data_33, 
         nvm_data_32, nvm_data_31, nvm_data_30, nvm_data_29, nvm_data_28, 
         nvm_data_27, nvm_data_26, nvm_data_25, nvm_data_24, nvm_data_23, 
         nvm_data_22, nvm_data_21, nvm_data_20, nvm_data_19, nvm_data_18, 
         nvm_data_17, nvm_data_16, nvm_data_15, nvm_data_14, nvm_data_13, 
         nvm_data_12, nvm_data_11, nvm_data_10, nvm_data_9, nvm_data_8, 
         nvm_data_7, nvm_data_6, nvm_data_5, nvm_data_4, nvm_data_3, nvm_data_2, 
         nvm_data_1, nvm_data_0, nvm_module_GND0, 
         camera_module_algo_module_prev_cont_enable, nx879, 
         camera_module_algo_module_modCU_current_state_13, 
         camera_module_algo_module_address_value_1, 
         camera_module_algo_module_modCU_current_state_10, 
         camera_module_algo_module_modCU_current_state_7, 
         camera_module_algo_module_modCU_current_state_6, 
         camera_module_algo_module_modCU_current_state_5, 
         camera_module_algo_module_pixel_enable, 
         camera_module_algo_module_modCU_current_state_12, 
         camera_module_algo_module_nvm_address_enable, nx883, 
         camera_module_ack_from_DMA, camera_module_cache_address_from_DMA_7, 
         camera_module_write_from_DMA, camera_module_DMA_module_signals_4, 
         camera_module_DMA_module_controlUnit_state_1, 
         camera_module_DMA_module_signals_1, nx20, nx36, nx48, 
         camera_module_cache_address_from_DMA_0, nx56, nx78, nx889, nx80, nx126, 
         nx128, nx130, camera_module_DMA_module_controlUnit_state_4, nx160, 
         nx178, camera_module_cache_address_from_DMA_4, nx216, 
         camera_module_cache_address_from_DMA_5, nx897, nx218, nx226, 
         camera_module_cache_address_from_DMA_6, nx264, nx268, nx276, nx294, 
         nx308, nx348, camera_module_algo_module_regs_rst, nx404, nx408, 
         camera_module_algo_module_address_value_0, nx418, nx426, nx436, nx448, 
         camera_module_algo_module_address_value_3, nx460, 
         camera_module_algo_module_address_value_2, nx903, nx462, nx470, nx496, 
         nx512, camera_module_algo_module_address_value_7, nx518, 
         camera_module_algo_module_address_value_4, nx905, nx520, nx528, 
         camera_module_algo_module_address_value_5, nx552, nx566, 
         camera_module_algo_module_address_value_6, nx908, nx568, nx576, nx602, 
         nx622, camera_module_algo_module_current_cont_value_15, 
         camera_module_algo_module_Addout_value_15, 
         camera_module_algo_module_current_cont_value_0, 
         camera_module_algo_module_Addout_value_0, nx656, nx664, nx678, 
         camera_module_algo_module_diff_value_0, nx686, nx688, 
         camera_module_algo_module_pixel_value_8, nx704, 
         camera_module_algo_module_pixel_value_0, nx738, nx752, nx770, nx802, 
         nx810, nx828, nx836, nx842, nx860, nx872, nx880, nx888, nx894, nx898, 
         nx906, nx912, camera_module_cache_ram_255__0, nx932, nx934, nx946, 
         nx954, nx962, nx968, nx972, nx980, nx986, nx1004, nx1016, nx1024, 
         nx1032, nx1038, nx1042, nx1050, nx1056, nx1088, nx1098, nx1110, nx1114, 
         nx1120, nx1130, nx1142, nx1146, nx1158, nx1170, nx1174, nx1186, 
         camera_module_cache_ram_239__0, camera_module_cache_ram_223__0, 
         camera_module_cache_ram_207__0, camera_module_cache_ram_191__0, nx1270, 
         camera_module_cache_ram_175__0, nx1288, camera_module_cache_ram_159__0, 
         nx1308, camera_module_cache_ram_143__0, nx1326, nx1348, 
         camera_module_cache_ram_127__0, nx1354, camera_module_cache_ram_111__0, 
         nx1372, camera_module_cache_ram_95__0, nx1392, 
         camera_module_cache_ram_79__0, nx1410, camera_module_cache_ram_63__0, 
         nx1434, camera_module_cache_ram_47__0, nx1452, 
         camera_module_cache_ram_31__0, nx1472, camera_module_cache_ram_15__0, 
         nx1490, nx1512, camera_module_cache_ram_254__0, 
         camera_module_cache_ram_238__0, camera_module_cache_ram_222__0, 
         camera_module_cache_ram_206__0, camera_module_cache_ram_190__0, 
         camera_module_cache_ram_174__0, camera_module_cache_ram_158__0, 
         camera_module_cache_ram_142__0, nx1666, camera_module_cache_ram_126__0, 
         camera_module_cache_ram_110__0, camera_module_cache_ram_94__0, 
         camera_module_cache_ram_78__0, camera_module_cache_ram_62__0, 
         camera_module_cache_ram_46__0, camera_module_cache_ram_30__0, 
         camera_module_cache_ram_14__0, nx1808, camera_module_cache_ram_253__0, 
         camera_module_cache_ram_237__0, camera_module_cache_ram_221__0, 
         camera_module_cache_ram_205__0, camera_module_cache_ram_189__0, 
         camera_module_cache_ram_173__0, camera_module_cache_ram_157__0, 
         camera_module_cache_ram_141__0, nx1964, camera_module_cache_ram_125__0, 
         camera_module_cache_ram_109__0, camera_module_cache_ram_93__0, 
         camera_module_cache_ram_77__0, camera_module_cache_ram_61__0, 
         camera_module_cache_ram_45__0, camera_module_cache_ram_29__0, 
         camera_module_cache_ram_13__0, nx2106, camera_module_cache_ram_252__0, 
         camera_module_cache_ram_236__0, camera_module_cache_ram_220__0, 
         camera_module_cache_ram_204__0, camera_module_cache_ram_188__0, 
         camera_module_cache_ram_172__0, camera_module_cache_ram_156__0, 
         camera_module_cache_ram_140__0, nx2258, camera_module_cache_ram_124__0, 
         camera_module_cache_ram_108__0, camera_module_cache_ram_92__0, 
         camera_module_cache_ram_76__0, camera_module_cache_ram_60__0, 
         camera_module_cache_ram_44__0, camera_module_cache_ram_28__0, 
         camera_module_cache_ram_12__0, nx2400, nx2410, nx2416, 
         camera_module_cache_ram_251__0, nx2424, camera_module_cache_ram_235__0, 
         nx2440, camera_module_cache_ram_219__0, nx2458, 
         camera_module_cache_ram_203__0, nx2474, camera_module_cache_ram_187__0, 
         nx2494, camera_module_cache_ram_171__0, nx2510, 
         camera_module_cache_ram_155__0, nx2528, camera_module_cache_ram_139__0, 
         nx2544, nx2558, camera_module_cache_ram_123__0, nx2566, 
         camera_module_cache_ram_107__0, nx2582, camera_module_cache_ram_91__0, 
         nx2600, camera_module_cache_ram_75__0, nx2616, 
         camera_module_cache_ram_59__0, nx2636, camera_module_cache_ram_43__0, 
         nx2652, camera_module_cache_ram_27__0, nx2670, 
         camera_module_cache_ram_11__0, nx2686, nx2700, nx2708, 
         camera_module_cache_ram_250__0, nx2716, camera_module_cache_ram_234__0, 
         nx2732, camera_module_cache_ram_218__0, nx2750, 
         camera_module_cache_ram_202__0, nx2766, camera_module_cache_ram_186__0, 
         nx2786, camera_module_cache_ram_170__0, nx2802, 
         camera_module_cache_ram_154__0, nx2820, camera_module_cache_ram_138__0, 
         nx2836, nx2850, camera_module_cache_ram_122__0, nx2858, 
         camera_module_cache_ram_106__0, nx2874, camera_module_cache_ram_90__0, 
         nx2892, camera_module_cache_ram_74__0, nx2908, 
         camera_module_cache_ram_58__0, nx2928, camera_module_cache_ram_42__0, 
         nx2944, camera_module_cache_ram_26__0, nx2962, 
         camera_module_cache_ram_10__0, nx2978, nx2992, nx3002, 
         camera_module_cache_ram_249__0, nx3010, camera_module_cache_ram_233__0, 
         nx3026, camera_module_cache_ram_217__0, nx3044, 
         camera_module_cache_ram_201__0, nx3060, camera_module_cache_ram_185__0, 
         nx3080, camera_module_cache_ram_169__0, nx3096, 
         camera_module_cache_ram_153__0, nx3114, camera_module_cache_ram_137__0, 
         nx3130, nx3144, camera_module_cache_ram_121__0, nx3152, 
         camera_module_cache_ram_105__0, nx3168, camera_module_cache_ram_89__0, 
         nx3186, camera_module_cache_ram_73__0, nx3202, 
         camera_module_cache_ram_57__0, nx3222, camera_module_cache_ram_41__0, 
         nx3238, camera_module_cache_ram_25__0, nx3256, 
         camera_module_cache_ram_9__0, nx3272, nx3286, nx3294, 
         camera_module_cache_ram_248__0, nx3302, camera_module_cache_ram_232__0, 
         nx3318, camera_module_cache_ram_216__0, nx3336, 
         camera_module_cache_ram_200__0, nx3352, camera_module_cache_ram_184__0, 
         nx3372, camera_module_cache_ram_168__0, nx3388, 
         camera_module_cache_ram_152__0, nx3406, camera_module_cache_ram_136__0, 
         nx3422, nx3436, camera_module_cache_ram_120__0, nx3444, 
         camera_module_cache_ram_104__0, nx3460, camera_module_cache_ram_88__0, 
         nx3478, camera_module_cache_ram_72__0, nx3494, 
         camera_module_cache_ram_56__0, nx3514, camera_module_cache_ram_40__0, 
         nx3530, camera_module_cache_ram_24__0, nx3548, 
         camera_module_cache_ram_8__0, nx3564, nx3578, nx3588, nx3596, 
         camera_module_cache_ram_247__0, nx3604, camera_module_cache_ram_231__0, 
         nx3620, camera_module_cache_ram_215__0, nx3638, 
         camera_module_cache_ram_199__0, nx3654, camera_module_cache_ram_183__0, 
         nx3674, camera_module_cache_ram_167__0, nx3690, 
         camera_module_cache_ram_151__0, nx3708, camera_module_cache_ram_135__0, 
         nx3724, nx3738, camera_module_cache_ram_119__0, nx3746, 
         camera_module_cache_ram_103__0, nx3762, camera_module_cache_ram_87__0, 
         nx3780, camera_module_cache_ram_71__0, nx3796, 
         camera_module_cache_ram_55__0, nx3816, camera_module_cache_ram_39__0, 
         nx3832, camera_module_cache_ram_23__0, nx3850, 
         camera_module_cache_ram_7__0, nx3866, nx3880, nx3888, 
         camera_module_cache_ram_246__0, nx3896, camera_module_cache_ram_230__0, 
         nx3912, camera_module_cache_ram_214__0, nx3930, 
         camera_module_cache_ram_198__0, nx3946, camera_module_cache_ram_182__0, 
         nx3966, camera_module_cache_ram_166__0, nx3982, 
         camera_module_cache_ram_150__0, nx4000, camera_module_cache_ram_134__0, 
         nx4016, nx4030, camera_module_cache_ram_118__0, nx4038, 
         camera_module_cache_ram_102__0, nx4054, camera_module_cache_ram_86__0, 
         nx4072, camera_module_cache_ram_70__0, nx4088, 
         camera_module_cache_ram_54__0, nx4108, camera_module_cache_ram_38__0, 
         nx4124, camera_module_cache_ram_22__0, nx4142, 
         camera_module_cache_ram_6__0, nx4158, nx4172, nx4182, 
         camera_module_cache_ram_245__0, nx4190, camera_module_cache_ram_229__0, 
         nx4206, camera_module_cache_ram_213__0, nx4224, 
         camera_module_cache_ram_197__0, nx4240, camera_module_cache_ram_181__0, 
         nx4260, camera_module_cache_ram_165__0, nx4276, 
         camera_module_cache_ram_149__0, nx4294, camera_module_cache_ram_133__0, 
         nx4310, nx4324, camera_module_cache_ram_117__0, nx4332, 
         camera_module_cache_ram_101__0, nx4348, camera_module_cache_ram_85__0, 
         nx4366, camera_module_cache_ram_69__0, nx4382, 
         camera_module_cache_ram_53__0, nx4402, camera_module_cache_ram_37__0, 
         nx4418, camera_module_cache_ram_21__0, nx4436, 
         camera_module_cache_ram_5__0, nx4452, nx4466, nx4474, 
         camera_module_cache_ram_244__0, nx4482, camera_module_cache_ram_228__0, 
         nx4498, camera_module_cache_ram_212__0, nx4516, 
         camera_module_cache_ram_196__0, nx4532, camera_module_cache_ram_180__0, 
         nx4552, camera_module_cache_ram_164__0, nx4568, 
         camera_module_cache_ram_148__0, nx4586, camera_module_cache_ram_132__0, 
         nx4602, nx4616, camera_module_cache_ram_116__0, nx4624, 
         camera_module_cache_ram_100__0, nx4640, camera_module_cache_ram_84__0, 
         nx4658, camera_module_cache_ram_68__0, nx4674, 
         camera_module_cache_ram_52__0, nx4694, camera_module_cache_ram_36__0, 
         nx4710, camera_module_cache_ram_20__0, nx4728, 
         camera_module_cache_ram_4__0, nx4744, nx4758, nx4768, nx4772, 
         camera_module_cache_ram_243__0, nx4780, camera_module_cache_ram_227__0, 
         nx4796, camera_module_cache_ram_211__0, nx4814, 
         camera_module_cache_ram_195__0, nx4830, camera_module_cache_ram_179__0, 
         nx4850, camera_module_cache_ram_163__0, nx4866, 
         camera_module_cache_ram_147__0, nx4884, camera_module_cache_ram_131__0, 
         nx4900, nx4914, camera_module_cache_ram_115__0, nx4922, 
         camera_module_cache_ram_99__0, nx4938, camera_module_cache_ram_83__0, 
         nx4956, camera_module_cache_ram_67__0, nx4972, 
         camera_module_cache_ram_51__0, nx4992, camera_module_cache_ram_35__0, 
         nx5008, camera_module_cache_ram_19__0, nx5026, 
         camera_module_cache_ram_3__0, nx5042, nx5056, nx5064, 
         camera_module_cache_ram_242__0, nx5072, camera_module_cache_ram_226__0, 
         nx5088, camera_module_cache_ram_210__0, nx5106, 
         camera_module_cache_ram_194__0, nx5122, camera_module_cache_ram_178__0, 
         nx5142, camera_module_cache_ram_162__0, nx5158, 
         camera_module_cache_ram_146__0, nx5176, camera_module_cache_ram_130__0, 
         nx5192, nx5206, camera_module_cache_ram_114__0, nx5214, 
         camera_module_cache_ram_98__0, nx5230, camera_module_cache_ram_82__0, 
         nx5248, camera_module_cache_ram_66__0, nx5264, 
         camera_module_cache_ram_50__0, nx5284, camera_module_cache_ram_34__0, 
         nx5300, camera_module_cache_ram_18__0, nx5318, 
         camera_module_cache_ram_2__0, nx5334, nx5348, nx5358, 
         camera_module_cache_ram_241__0, nx5366, camera_module_cache_ram_225__0, 
         nx5382, camera_module_cache_ram_209__0, nx5400, 
         camera_module_cache_ram_193__0, nx5416, camera_module_cache_ram_177__0, 
         nx5436, camera_module_cache_ram_161__0, nx5452, 
         camera_module_cache_ram_145__0, nx5470, camera_module_cache_ram_129__0, 
         nx5486, nx5500, camera_module_cache_ram_113__0, nx5508, 
         camera_module_cache_ram_97__0, nx5524, camera_module_cache_ram_81__0, 
         nx5542, camera_module_cache_ram_65__0, nx5558, 
         camera_module_cache_ram_49__0, nx5578, camera_module_cache_ram_33__0, 
         nx5594, camera_module_cache_ram_17__0, nx5612, 
         camera_module_cache_ram_1__0, nx5628, nx5642, nx5650, 
         camera_module_cache_ram_240__0, nx5658, camera_module_cache_ram_224__0, 
         nx5674, camera_module_cache_ram_208__0, nx5692, 
         camera_module_cache_ram_192__0, nx5708, camera_module_cache_ram_176__0, 
         nx5728, camera_module_cache_ram_160__0, nx5744, 
         camera_module_cache_ram_144__0, nx5762, camera_module_cache_ram_128__0, 
         nx5778, nx5792, camera_module_cache_ram_112__0, nx5800, 
         camera_module_cache_ram_96__0, nx5816, camera_module_cache_ram_80__0, 
         nx5834, camera_module_cache_ram_64__0, nx5850, 
         camera_module_cache_ram_48__0, nx5870, camera_module_cache_ram_32__0, 
         nx5886, camera_module_cache_ram_16__0, nx5904, 
         camera_module_cache_ram_0__0, nx5920, nx5934, nx5944, nx5964, nx5972, 
         camera_module_algo_module_pixel_value_1, camera_module_cache_ram_255__1, 
         nx6002, nx6012, nx6024, nx6028, nx6034, nx6044, nx6056, nx6060, nx6072, 
         nx6084, nx6088, nx6100, camera_module_cache_ram_239__1, 
         camera_module_cache_ram_223__1, camera_module_cache_ram_207__1, 
         camera_module_cache_ram_191__1, camera_module_cache_ram_175__1, 
         camera_module_cache_ram_159__1, camera_module_cache_ram_143__1, nx6178, 
         camera_module_cache_ram_127__1, camera_module_cache_ram_111__1, 
         camera_module_cache_ram_95__1, camera_module_cache_ram_79__1, 
         camera_module_cache_ram_63__1, camera_module_cache_ram_47__1, 
         camera_module_cache_ram_31__1, camera_module_cache_ram_15__1, nx6256, 
         camera_module_cache_ram_254__1, camera_module_cache_ram_238__1, 
         camera_module_cache_ram_222__1, camera_module_cache_ram_206__1, 
         camera_module_cache_ram_190__1, camera_module_cache_ram_174__1, 
         camera_module_cache_ram_158__1, camera_module_cache_ram_142__1, nx6340, 
         camera_module_cache_ram_126__1, camera_module_cache_ram_110__1, 
         camera_module_cache_ram_94__1, camera_module_cache_ram_78__1, 
         camera_module_cache_ram_62__1, camera_module_cache_ram_46__1, 
         camera_module_cache_ram_30__1, camera_module_cache_ram_14__1, nx6418, 
         camera_module_cache_ram_253__1, camera_module_cache_ram_237__1, 
         camera_module_cache_ram_221__1, camera_module_cache_ram_205__1, 
         camera_module_cache_ram_189__1, camera_module_cache_ram_173__1, 
         camera_module_cache_ram_157__1, camera_module_cache_ram_141__1, nx6504, 
         camera_module_cache_ram_125__1, camera_module_cache_ram_109__1, 
         camera_module_cache_ram_93__1, camera_module_cache_ram_77__1, 
         camera_module_cache_ram_61__1, camera_module_cache_ram_45__1, 
         camera_module_cache_ram_29__1, camera_module_cache_ram_13__1, nx6582, 
         camera_module_cache_ram_252__1, camera_module_cache_ram_236__1, 
         camera_module_cache_ram_220__1, camera_module_cache_ram_204__1, 
         camera_module_cache_ram_188__1, camera_module_cache_ram_172__1, 
         camera_module_cache_ram_156__1, camera_module_cache_ram_140__1, nx6666, 
         camera_module_cache_ram_124__1, camera_module_cache_ram_108__1, 
         camera_module_cache_ram_92__1, camera_module_cache_ram_76__1, 
         camera_module_cache_ram_60__1, camera_module_cache_ram_44__1, 
         camera_module_cache_ram_28__1, camera_module_cache_ram_12__1, nx6744, 
         nx6754, camera_module_cache_ram_251__1, camera_module_cache_ram_235__1, 
         camera_module_cache_ram_219__1, camera_module_cache_ram_203__1, 
         camera_module_cache_ram_187__1, camera_module_cache_ram_171__1, 
         camera_module_cache_ram_155__1, camera_module_cache_ram_139__1, nx6832, 
         camera_module_cache_ram_123__1, camera_module_cache_ram_107__1, 
         camera_module_cache_ram_91__1, camera_module_cache_ram_75__1, 
         camera_module_cache_ram_59__1, camera_module_cache_ram_43__1, 
         camera_module_cache_ram_27__1, camera_module_cache_ram_11__1, nx6910, 
         camera_module_cache_ram_250__1, camera_module_cache_ram_234__1, 
         camera_module_cache_ram_218__1, camera_module_cache_ram_202__1, 
         camera_module_cache_ram_186__1, camera_module_cache_ram_170__1, 
         camera_module_cache_ram_154__1, camera_module_cache_ram_138__1, nx6994, 
         camera_module_cache_ram_122__1, camera_module_cache_ram_106__1, 
         camera_module_cache_ram_90__1, camera_module_cache_ram_74__1, 
         camera_module_cache_ram_58__1, camera_module_cache_ram_42__1, 
         camera_module_cache_ram_26__1, camera_module_cache_ram_10__1, nx7072, 
         camera_module_cache_ram_249__1, camera_module_cache_ram_233__1, 
         camera_module_cache_ram_217__1, camera_module_cache_ram_201__1, 
         camera_module_cache_ram_185__1, camera_module_cache_ram_169__1, 
         camera_module_cache_ram_153__1, camera_module_cache_ram_137__1, nx7158, 
         camera_module_cache_ram_121__1, camera_module_cache_ram_105__1, 
         camera_module_cache_ram_89__1, camera_module_cache_ram_73__1, 
         camera_module_cache_ram_57__1, camera_module_cache_ram_41__1, 
         camera_module_cache_ram_25__1, camera_module_cache_ram_9__1, nx7236, 
         camera_module_cache_ram_248__1, camera_module_cache_ram_232__1, 
         camera_module_cache_ram_216__1, camera_module_cache_ram_200__1, 
         camera_module_cache_ram_184__1, camera_module_cache_ram_168__1, 
         camera_module_cache_ram_152__1, camera_module_cache_ram_136__1, nx7320, 
         camera_module_cache_ram_120__1, camera_module_cache_ram_104__1, 
         camera_module_cache_ram_88__1, camera_module_cache_ram_72__1, 
         camera_module_cache_ram_56__1, camera_module_cache_ram_40__1, 
         camera_module_cache_ram_24__1, camera_module_cache_ram_8__1, nx7398, 
         nx7408, camera_module_cache_ram_247__1, camera_module_cache_ram_231__1, 
         camera_module_cache_ram_215__1, camera_module_cache_ram_199__1, 
         camera_module_cache_ram_183__1, camera_module_cache_ram_167__1, 
         camera_module_cache_ram_151__1, camera_module_cache_ram_135__1, nx7488, 
         camera_module_cache_ram_119__1, camera_module_cache_ram_103__1, 
         camera_module_cache_ram_87__1, camera_module_cache_ram_71__1, 
         camera_module_cache_ram_55__1, camera_module_cache_ram_39__1, 
         camera_module_cache_ram_23__1, camera_module_cache_ram_7__1, nx7566, 
         camera_module_cache_ram_246__1, camera_module_cache_ram_230__1, 
         camera_module_cache_ram_214__1, camera_module_cache_ram_198__1, 
         camera_module_cache_ram_182__1, camera_module_cache_ram_166__1, 
         camera_module_cache_ram_150__1, camera_module_cache_ram_134__1, nx7650, 
         camera_module_cache_ram_118__1, camera_module_cache_ram_102__1, 
         camera_module_cache_ram_86__1, camera_module_cache_ram_70__1, 
         camera_module_cache_ram_54__1, camera_module_cache_ram_38__1, 
         camera_module_cache_ram_22__1, camera_module_cache_ram_6__1, nx7728, 
         camera_module_cache_ram_245__1, camera_module_cache_ram_229__1, 
         camera_module_cache_ram_213__1, camera_module_cache_ram_197__1, 
         camera_module_cache_ram_181__1, camera_module_cache_ram_165__1, 
         camera_module_cache_ram_149__1, camera_module_cache_ram_133__1, nx7814, 
         camera_module_cache_ram_117__1, camera_module_cache_ram_101__1, 
         camera_module_cache_ram_85__1, camera_module_cache_ram_69__1, 
         camera_module_cache_ram_53__1, camera_module_cache_ram_37__1, 
         camera_module_cache_ram_21__1, camera_module_cache_ram_5__1, nx7892, 
         camera_module_cache_ram_244__1, camera_module_cache_ram_228__1, 
         camera_module_cache_ram_212__1, camera_module_cache_ram_196__1, 
         camera_module_cache_ram_180__1, camera_module_cache_ram_164__1, 
         camera_module_cache_ram_148__1, camera_module_cache_ram_132__1, nx7976, 
         camera_module_cache_ram_116__1, camera_module_cache_ram_100__1, 
         camera_module_cache_ram_84__1, camera_module_cache_ram_68__1, 
         camera_module_cache_ram_52__1, camera_module_cache_ram_36__1, 
         camera_module_cache_ram_20__1, camera_module_cache_ram_4__1, nx8054, 
         nx8064, camera_module_cache_ram_243__1, camera_module_cache_ram_227__1, 
         camera_module_cache_ram_211__1, camera_module_cache_ram_195__1, 
         camera_module_cache_ram_179__1, camera_module_cache_ram_163__1, 
         camera_module_cache_ram_147__1, camera_module_cache_ram_131__1, nx8142, 
         camera_module_cache_ram_115__1, camera_module_cache_ram_99__1, 
         camera_module_cache_ram_83__1, camera_module_cache_ram_67__1, 
         camera_module_cache_ram_51__1, camera_module_cache_ram_35__1, 
         camera_module_cache_ram_19__1, camera_module_cache_ram_3__1, nx8220, 
         camera_module_cache_ram_242__1, camera_module_cache_ram_226__1, 
         camera_module_cache_ram_210__1, camera_module_cache_ram_194__1, 
         camera_module_cache_ram_178__1, camera_module_cache_ram_162__1, 
         camera_module_cache_ram_146__1, camera_module_cache_ram_130__1, nx8304, 
         camera_module_cache_ram_114__1, camera_module_cache_ram_98__1, 
         camera_module_cache_ram_82__1, camera_module_cache_ram_66__1, 
         camera_module_cache_ram_50__1, camera_module_cache_ram_34__1, 
         camera_module_cache_ram_18__1, camera_module_cache_ram_2__1, nx8382, 
         camera_module_cache_ram_241__1, camera_module_cache_ram_225__1, 
         camera_module_cache_ram_209__1, camera_module_cache_ram_193__1, 
         camera_module_cache_ram_177__1, camera_module_cache_ram_161__1, 
         camera_module_cache_ram_145__1, camera_module_cache_ram_129__1, nx8468, 
         camera_module_cache_ram_113__1, camera_module_cache_ram_97__1, 
         camera_module_cache_ram_81__1, camera_module_cache_ram_65__1, 
         camera_module_cache_ram_49__1, camera_module_cache_ram_33__1, 
         camera_module_cache_ram_17__1, camera_module_cache_ram_1__1, nx8546, 
         camera_module_cache_ram_240__1, camera_module_cache_ram_224__1, 
         camera_module_cache_ram_208__1, camera_module_cache_ram_192__1, 
         camera_module_cache_ram_176__1, camera_module_cache_ram_160__1, 
         camera_module_cache_ram_144__1, camera_module_cache_ram_128__1, nx8630, 
         camera_module_cache_ram_112__1, camera_module_cache_ram_96__1, 
         camera_module_cache_ram_80__1, camera_module_cache_ram_64__1, 
         camera_module_cache_ram_48__1, camera_module_cache_ram_32__1, 
         camera_module_cache_ram_16__1, camera_module_cache_ram_0__1, nx8708, 
         nx8718, nx8730, nx8738, nx8754, camera_module_algo_module_pixel_value_2, 
         camera_module_cache_ram_255__2, nx8776, nx8786, nx8798, nx8802, nx8808, 
         nx8818, nx8830, nx8834, nx8846, nx8858, nx8862, nx8874, 
         camera_module_cache_ram_239__2, camera_module_cache_ram_223__2, 
         camera_module_cache_ram_207__2, camera_module_cache_ram_191__2, 
         camera_module_cache_ram_175__2, camera_module_cache_ram_159__2, 
         camera_module_cache_ram_143__2, nx8952, camera_module_cache_ram_127__2, 
         camera_module_cache_ram_111__2, camera_module_cache_ram_95__2, 
         camera_module_cache_ram_79__2, camera_module_cache_ram_63__2, 
         camera_module_cache_ram_47__2, camera_module_cache_ram_31__2, 
         camera_module_cache_ram_15__2, nx9030, camera_module_cache_ram_254__2, 
         camera_module_cache_ram_238__2, camera_module_cache_ram_222__2, 
         camera_module_cache_ram_206__2, camera_module_cache_ram_190__2, 
         camera_module_cache_ram_174__2, camera_module_cache_ram_158__2, 
         camera_module_cache_ram_142__2, nx9114, camera_module_cache_ram_126__2, 
         camera_module_cache_ram_110__2, camera_module_cache_ram_94__2, 
         camera_module_cache_ram_78__2, camera_module_cache_ram_62__2, 
         camera_module_cache_ram_46__2, camera_module_cache_ram_30__2, 
         camera_module_cache_ram_14__2, nx9192, camera_module_cache_ram_253__2, 
         camera_module_cache_ram_237__2, camera_module_cache_ram_221__2, 
         camera_module_cache_ram_205__2, camera_module_cache_ram_189__2, 
         camera_module_cache_ram_173__2, camera_module_cache_ram_157__2, 
         camera_module_cache_ram_141__2, nx9278, camera_module_cache_ram_125__2, 
         camera_module_cache_ram_109__2, camera_module_cache_ram_93__2, 
         camera_module_cache_ram_77__2, camera_module_cache_ram_61__2, 
         camera_module_cache_ram_45__2, camera_module_cache_ram_29__2, 
         camera_module_cache_ram_13__2, nx9356, camera_module_cache_ram_252__2, 
         camera_module_cache_ram_236__2, camera_module_cache_ram_220__2, 
         camera_module_cache_ram_204__2, camera_module_cache_ram_188__2, 
         camera_module_cache_ram_172__2, camera_module_cache_ram_156__2, 
         camera_module_cache_ram_140__2, nx9440, camera_module_cache_ram_124__2, 
         camera_module_cache_ram_108__2, camera_module_cache_ram_92__2, 
         camera_module_cache_ram_76__2, camera_module_cache_ram_60__2, 
         camera_module_cache_ram_44__2, camera_module_cache_ram_28__2, 
         camera_module_cache_ram_12__2, nx9518, nx9528, 
         camera_module_cache_ram_251__2, camera_module_cache_ram_235__2, 
         camera_module_cache_ram_219__2, camera_module_cache_ram_203__2, 
         camera_module_cache_ram_187__2, camera_module_cache_ram_171__2, 
         camera_module_cache_ram_155__2, camera_module_cache_ram_139__2, nx9606, 
         camera_module_cache_ram_123__2, camera_module_cache_ram_107__2, 
         camera_module_cache_ram_91__2, camera_module_cache_ram_75__2, 
         camera_module_cache_ram_59__2, camera_module_cache_ram_43__2, 
         camera_module_cache_ram_27__2, camera_module_cache_ram_11__2, nx9684, 
         camera_module_cache_ram_250__2, camera_module_cache_ram_234__2, 
         camera_module_cache_ram_218__2, camera_module_cache_ram_202__2, 
         camera_module_cache_ram_186__2, camera_module_cache_ram_170__2, 
         camera_module_cache_ram_154__2, camera_module_cache_ram_138__2, nx9768, 
         camera_module_cache_ram_122__2, camera_module_cache_ram_106__2, 
         camera_module_cache_ram_90__2, camera_module_cache_ram_74__2, 
         camera_module_cache_ram_58__2, camera_module_cache_ram_42__2, 
         camera_module_cache_ram_26__2, camera_module_cache_ram_10__2, nx9846, 
         camera_module_cache_ram_249__2, camera_module_cache_ram_233__2, 
         camera_module_cache_ram_217__2, camera_module_cache_ram_201__2, 
         camera_module_cache_ram_185__2, camera_module_cache_ram_169__2, 
         camera_module_cache_ram_153__2, camera_module_cache_ram_137__2, nx9932, 
         camera_module_cache_ram_121__2, camera_module_cache_ram_105__2, 
         camera_module_cache_ram_89__2, camera_module_cache_ram_73__2, 
         camera_module_cache_ram_57__2, camera_module_cache_ram_41__2, 
         camera_module_cache_ram_25__2, camera_module_cache_ram_9__2, nx10010, 
         camera_module_cache_ram_248__2, camera_module_cache_ram_232__2, 
         camera_module_cache_ram_216__2, camera_module_cache_ram_200__2, 
         camera_module_cache_ram_184__2, camera_module_cache_ram_168__2, 
         camera_module_cache_ram_152__2, camera_module_cache_ram_136__2, nx10094, 
         camera_module_cache_ram_120__2, camera_module_cache_ram_104__2, 
         camera_module_cache_ram_88__2, camera_module_cache_ram_72__2, 
         camera_module_cache_ram_56__2, camera_module_cache_ram_40__2, 
         camera_module_cache_ram_24__2, camera_module_cache_ram_8__2, nx10172, 
         nx10182, camera_module_cache_ram_247__2, camera_module_cache_ram_231__2, 
         camera_module_cache_ram_215__2, camera_module_cache_ram_199__2, 
         camera_module_cache_ram_183__2, camera_module_cache_ram_167__2, 
         camera_module_cache_ram_151__2, camera_module_cache_ram_135__2, nx10262, 
         camera_module_cache_ram_119__2, camera_module_cache_ram_103__2, 
         camera_module_cache_ram_87__2, camera_module_cache_ram_71__2, 
         camera_module_cache_ram_55__2, camera_module_cache_ram_39__2, 
         camera_module_cache_ram_23__2, camera_module_cache_ram_7__2, nx10340, 
         camera_module_cache_ram_246__2, camera_module_cache_ram_230__2, 
         camera_module_cache_ram_214__2, camera_module_cache_ram_198__2, 
         camera_module_cache_ram_182__2, camera_module_cache_ram_166__2, 
         camera_module_cache_ram_150__2, camera_module_cache_ram_134__2, nx10424, 
         camera_module_cache_ram_118__2, camera_module_cache_ram_102__2, 
         camera_module_cache_ram_86__2, camera_module_cache_ram_70__2, 
         camera_module_cache_ram_54__2, camera_module_cache_ram_38__2, 
         camera_module_cache_ram_22__2, camera_module_cache_ram_6__2, nx10502, 
         camera_module_cache_ram_245__2, camera_module_cache_ram_229__2, 
         camera_module_cache_ram_213__2, camera_module_cache_ram_197__2, 
         camera_module_cache_ram_181__2, camera_module_cache_ram_165__2, 
         camera_module_cache_ram_149__2, camera_module_cache_ram_133__2, nx10588, 
         camera_module_cache_ram_117__2, camera_module_cache_ram_101__2, 
         camera_module_cache_ram_85__2, camera_module_cache_ram_69__2, 
         camera_module_cache_ram_53__2, camera_module_cache_ram_37__2, 
         camera_module_cache_ram_21__2, camera_module_cache_ram_5__2, nx10666, 
         camera_module_cache_ram_244__2, camera_module_cache_ram_228__2, 
         camera_module_cache_ram_212__2, camera_module_cache_ram_196__2, 
         camera_module_cache_ram_180__2, camera_module_cache_ram_164__2, 
         camera_module_cache_ram_148__2, camera_module_cache_ram_132__2, nx10750, 
         camera_module_cache_ram_116__2, camera_module_cache_ram_100__2, 
         camera_module_cache_ram_84__2, camera_module_cache_ram_68__2, 
         camera_module_cache_ram_52__2, camera_module_cache_ram_36__2, 
         camera_module_cache_ram_20__2, camera_module_cache_ram_4__2, nx10828, 
         nx10838, camera_module_cache_ram_243__2, camera_module_cache_ram_227__2, 
         camera_module_cache_ram_211__2, camera_module_cache_ram_195__2, 
         camera_module_cache_ram_179__2, camera_module_cache_ram_163__2, 
         camera_module_cache_ram_147__2, camera_module_cache_ram_131__2, nx10916, 
         camera_module_cache_ram_115__2, camera_module_cache_ram_99__2, 
         camera_module_cache_ram_83__2, camera_module_cache_ram_67__2, 
         camera_module_cache_ram_51__2, camera_module_cache_ram_35__2, 
         camera_module_cache_ram_19__2, camera_module_cache_ram_3__2, nx10994, 
         camera_module_cache_ram_242__2, camera_module_cache_ram_226__2, 
         camera_module_cache_ram_210__2, camera_module_cache_ram_194__2, 
         camera_module_cache_ram_178__2, camera_module_cache_ram_162__2, 
         camera_module_cache_ram_146__2, camera_module_cache_ram_130__2, nx11078, 
         camera_module_cache_ram_114__2, camera_module_cache_ram_98__2, 
         camera_module_cache_ram_82__2, camera_module_cache_ram_66__2, 
         camera_module_cache_ram_50__2, camera_module_cache_ram_34__2, 
         camera_module_cache_ram_18__2, camera_module_cache_ram_2__2, nx11156, 
         camera_module_cache_ram_241__2, camera_module_cache_ram_225__2, 
         camera_module_cache_ram_209__2, camera_module_cache_ram_193__2, 
         camera_module_cache_ram_177__2, camera_module_cache_ram_161__2, 
         camera_module_cache_ram_145__2, camera_module_cache_ram_129__2, nx11242, 
         camera_module_cache_ram_113__2, camera_module_cache_ram_97__2, 
         camera_module_cache_ram_81__2, camera_module_cache_ram_65__2, 
         camera_module_cache_ram_49__2, camera_module_cache_ram_33__2, 
         camera_module_cache_ram_17__2, camera_module_cache_ram_1__2, nx11320, 
         camera_module_cache_ram_240__2, camera_module_cache_ram_224__2, 
         camera_module_cache_ram_208__2, camera_module_cache_ram_192__2, 
         camera_module_cache_ram_176__2, camera_module_cache_ram_160__2, 
         camera_module_cache_ram_144__2, camera_module_cache_ram_128__2, nx11404, 
         camera_module_cache_ram_112__2, camera_module_cache_ram_96__2, 
         camera_module_cache_ram_80__2, camera_module_cache_ram_64__2, 
         camera_module_cache_ram_48__2, camera_module_cache_ram_32__2, 
         camera_module_cache_ram_16__2, camera_module_cache_ram_0__2, nx11482, 
         nx11492, nx11512, nx11520, camera_module_algo_module_pixel_value_3, 
         camera_module_cache_ram_255__3, nx11550, nx11560, nx11572, nx11576, 
         nx11582, nx11592, nx11604, nx11608, nx11620, nx11632, nx11636, nx11648, 
         camera_module_cache_ram_239__3, camera_module_cache_ram_223__3, 
         camera_module_cache_ram_207__3, camera_module_cache_ram_191__3, 
         camera_module_cache_ram_175__3, camera_module_cache_ram_159__3, 
         camera_module_cache_ram_143__3, nx11726, camera_module_cache_ram_127__3, 
         camera_module_cache_ram_111__3, camera_module_cache_ram_95__3, 
         camera_module_cache_ram_79__3, camera_module_cache_ram_63__3, 
         camera_module_cache_ram_47__3, camera_module_cache_ram_31__3, 
         camera_module_cache_ram_15__3, nx11804, camera_module_cache_ram_254__3, 
         camera_module_cache_ram_238__3, camera_module_cache_ram_222__3, 
         camera_module_cache_ram_206__3, camera_module_cache_ram_190__3, 
         camera_module_cache_ram_174__3, camera_module_cache_ram_158__3, 
         camera_module_cache_ram_142__3, nx11888, camera_module_cache_ram_126__3, 
         camera_module_cache_ram_110__3, camera_module_cache_ram_94__3, 
         camera_module_cache_ram_78__3, camera_module_cache_ram_62__3, 
         camera_module_cache_ram_46__3, camera_module_cache_ram_30__3, 
         camera_module_cache_ram_14__3, nx11966, camera_module_cache_ram_253__3, 
         camera_module_cache_ram_237__3, camera_module_cache_ram_221__3, 
         camera_module_cache_ram_205__3, camera_module_cache_ram_189__3, 
         camera_module_cache_ram_173__3, camera_module_cache_ram_157__3, 
         camera_module_cache_ram_141__3, nx12052, camera_module_cache_ram_125__3, 
         camera_module_cache_ram_109__3, camera_module_cache_ram_93__3, 
         camera_module_cache_ram_77__3, camera_module_cache_ram_61__3, 
         camera_module_cache_ram_45__3, camera_module_cache_ram_29__3, 
         camera_module_cache_ram_13__3, nx12130, camera_module_cache_ram_252__3, 
         camera_module_cache_ram_236__3, camera_module_cache_ram_220__3, 
         camera_module_cache_ram_204__3, camera_module_cache_ram_188__3, 
         camera_module_cache_ram_172__3, camera_module_cache_ram_156__3, 
         camera_module_cache_ram_140__3, nx12214, camera_module_cache_ram_124__3, 
         camera_module_cache_ram_108__3, camera_module_cache_ram_92__3, 
         camera_module_cache_ram_76__3, camera_module_cache_ram_60__3, 
         camera_module_cache_ram_44__3, camera_module_cache_ram_28__3, 
         camera_module_cache_ram_12__3, nx12292, nx12302, 
         camera_module_cache_ram_251__3, camera_module_cache_ram_235__3, 
         camera_module_cache_ram_219__3, camera_module_cache_ram_203__3, 
         camera_module_cache_ram_187__3, camera_module_cache_ram_171__3, 
         camera_module_cache_ram_155__3, camera_module_cache_ram_139__3, nx12380, 
         camera_module_cache_ram_123__3, camera_module_cache_ram_107__3, 
         camera_module_cache_ram_91__3, camera_module_cache_ram_75__3, 
         camera_module_cache_ram_59__3, camera_module_cache_ram_43__3, 
         camera_module_cache_ram_27__3, camera_module_cache_ram_11__3, nx12458, 
         camera_module_cache_ram_250__3, camera_module_cache_ram_234__3, 
         camera_module_cache_ram_218__3, camera_module_cache_ram_202__3, 
         camera_module_cache_ram_186__3, camera_module_cache_ram_170__3, 
         camera_module_cache_ram_154__3, camera_module_cache_ram_138__3, nx12542, 
         camera_module_cache_ram_122__3, camera_module_cache_ram_106__3, 
         camera_module_cache_ram_90__3, camera_module_cache_ram_74__3, 
         camera_module_cache_ram_58__3, camera_module_cache_ram_42__3, 
         camera_module_cache_ram_26__3, camera_module_cache_ram_10__3, nx12620, 
         camera_module_cache_ram_249__3, camera_module_cache_ram_233__3, 
         camera_module_cache_ram_217__3, camera_module_cache_ram_201__3, 
         camera_module_cache_ram_185__3, camera_module_cache_ram_169__3, 
         camera_module_cache_ram_153__3, camera_module_cache_ram_137__3, nx12706, 
         camera_module_cache_ram_121__3, camera_module_cache_ram_105__3, 
         camera_module_cache_ram_89__3, camera_module_cache_ram_73__3, 
         camera_module_cache_ram_57__3, camera_module_cache_ram_41__3, 
         camera_module_cache_ram_25__3, camera_module_cache_ram_9__3, nx12784, 
         camera_module_cache_ram_248__3, camera_module_cache_ram_232__3, 
         camera_module_cache_ram_216__3, camera_module_cache_ram_200__3, 
         camera_module_cache_ram_184__3, camera_module_cache_ram_168__3, 
         camera_module_cache_ram_152__3, camera_module_cache_ram_136__3, nx12868, 
         camera_module_cache_ram_120__3, camera_module_cache_ram_104__3, 
         camera_module_cache_ram_88__3, camera_module_cache_ram_72__3, 
         camera_module_cache_ram_56__3, camera_module_cache_ram_40__3, 
         camera_module_cache_ram_24__3, camera_module_cache_ram_8__3, nx12946, 
         nx12956, camera_module_cache_ram_247__3, camera_module_cache_ram_231__3, 
         camera_module_cache_ram_215__3, camera_module_cache_ram_199__3, 
         camera_module_cache_ram_183__3, camera_module_cache_ram_167__3, 
         camera_module_cache_ram_151__3, camera_module_cache_ram_135__3, nx13036, 
         camera_module_cache_ram_119__3, camera_module_cache_ram_103__3, 
         camera_module_cache_ram_87__3, camera_module_cache_ram_71__3, 
         camera_module_cache_ram_55__3, camera_module_cache_ram_39__3, 
         camera_module_cache_ram_23__3, camera_module_cache_ram_7__3, nx13114, 
         camera_module_cache_ram_246__3, camera_module_cache_ram_230__3, 
         camera_module_cache_ram_214__3, camera_module_cache_ram_198__3, 
         camera_module_cache_ram_182__3, camera_module_cache_ram_166__3, 
         camera_module_cache_ram_150__3, camera_module_cache_ram_134__3, nx13198, 
         camera_module_cache_ram_118__3, camera_module_cache_ram_102__3, 
         camera_module_cache_ram_86__3, camera_module_cache_ram_70__3, 
         camera_module_cache_ram_54__3, camera_module_cache_ram_38__3, 
         camera_module_cache_ram_22__3, camera_module_cache_ram_6__3, nx13276, 
         camera_module_cache_ram_245__3, camera_module_cache_ram_229__3, 
         camera_module_cache_ram_213__3, camera_module_cache_ram_197__3, 
         camera_module_cache_ram_181__3, camera_module_cache_ram_165__3, 
         camera_module_cache_ram_149__3, camera_module_cache_ram_133__3, nx13362, 
         camera_module_cache_ram_117__3, camera_module_cache_ram_101__3, 
         camera_module_cache_ram_85__3, camera_module_cache_ram_69__3, 
         camera_module_cache_ram_53__3, camera_module_cache_ram_37__3, 
         camera_module_cache_ram_21__3, camera_module_cache_ram_5__3, nx13440, 
         camera_module_cache_ram_244__3, camera_module_cache_ram_228__3, 
         camera_module_cache_ram_212__3, camera_module_cache_ram_196__3, 
         camera_module_cache_ram_180__3, camera_module_cache_ram_164__3, 
         camera_module_cache_ram_148__3, camera_module_cache_ram_132__3, nx13524, 
         camera_module_cache_ram_116__3, camera_module_cache_ram_100__3, 
         camera_module_cache_ram_84__3, camera_module_cache_ram_68__3, 
         camera_module_cache_ram_52__3, camera_module_cache_ram_36__3, 
         camera_module_cache_ram_20__3, camera_module_cache_ram_4__3, nx13602, 
         nx13612, camera_module_cache_ram_243__3, camera_module_cache_ram_227__3, 
         camera_module_cache_ram_211__3, camera_module_cache_ram_195__3, 
         camera_module_cache_ram_179__3, camera_module_cache_ram_163__3, 
         camera_module_cache_ram_147__3, camera_module_cache_ram_131__3, nx13690, 
         camera_module_cache_ram_115__3, camera_module_cache_ram_99__3, 
         camera_module_cache_ram_83__3, camera_module_cache_ram_67__3, 
         camera_module_cache_ram_51__3, camera_module_cache_ram_35__3, 
         camera_module_cache_ram_19__3, camera_module_cache_ram_3__3, nx13768, 
         camera_module_cache_ram_242__3, camera_module_cache_ram_226__3, 
         camera_module_cache_ram_210__3, camera_module_cache_ram_194__3, 
         camera_module_cache_ram_178__3, camera_module_cache_ram_162__3, 
         camera_module_cache_ram_146__3, camera_module_cache_ram_130__3, nx13852, 
         camera_module_cache_ram_114__3, camera_module_cache_ram_98__3, 
         camera_module_cache_ram_82__3, camera_module_cache_ram_66__3, 
         camera_module_cache_ram_50__3, camera_module_cache_ram_34__3, 
         camera_module_cache_ram_18__3, camera_module_cache_ram_2__3, nx13930, 
         camera_module_cache_ram_241__3, camera_module_cache_ram_225__3, 
         camera_module_cache_ram_209__3, camera_module_cache_ram_193__3, 
         camera_module_cache_ram_177__3, camera_module_cache_ram_161__3, 
         camera_module_cache_ram_145__3, camera_module_cache_ram_129__3, nx14016, 
         camera_module_cache_ram_113__3, camera_module_cache_ram_97__3, 
         camera_module_cache_ram_81__3, camera_module_cache_ram_65__3, 
         camera_module_cache_ram_49__3, camera_module_cache_ram_33__3, 
         camera_module_cache_ram_17__3, camera_module_cache_ram_1__3, nx14094, 
         camera_module_cache_ram_240__3, camera_module_cache_ram_224__3, 
         camera_module_cache_ram_208__3, camera_module_cache_ram_192__3, 
         camera_module_cache_ram_176__3, camera_module_cache_ram_160__3, 
         camera_module_cache_ram_144__3, camera_module_cache_ram_128__3, nx14178, 
         camera_module_cache_ram_112__3, camera_module_cache_ram_96__3, 
         camera_module_cache_ram_80__3, camera_module_cache_ram_64__3, 
         camera_module_cache_ram_48__3, camera_module_cache_ram_32__3, 
         camera_module_cache_ram_16__3, camera_module_cache_ram_0__3, nx14256, 
         nx14266, nx14278, nx14286, nx14302, 
         camera_module_algo_module_pixel_value_4, camera_module_cache_ram_255__4, 
         nx14324, nx14334, nx14346, nx14350, nx14356, nx14366, nx14378, nx14382, 
         nx14394, nx14406, nx14410, nx14422, camera_module_cache_ram_239__4, 
         camera_module_cache_ram_223__4, camera_module_cache_ram_207__4, 
         camera_module_cache_ram_191__4, camera_module_cache_ram_175__4, 
         camera_module_cache_ram_159__4, camera_module_cache_ram_143__4, nx14500, 
         camera_module_cache_ram_127__4, camera_module_cache_ram_111__4, 
         camera_module_cache_ram_95__4, camera_module_cache_ram_79__4, 
         camera_module_cache_ram_63__4, camera_module_cache_ram_47__4, 
         camera_module_cache_ram_31__4, camera_module_cache_ram_15__4, nx14578, 
         camera_module_cache_ram_254__4, camera_module_cache_ram_238__4, 
         camera_module_cache_ram_222__4, camera_module_cache_ram_206__4, 
         camera_module_cache_ram_190__4, camera_module_cache_ram_174__4, 
         camera_module_cache_ram_158__4, camera_module_cache_ram_142__4, nx14662, 
         camera_module_cache_ram_126__4, camera_module_cache_ram_110__4, 
         camera_module_cache_ram_94__4, camera_module_cache_ram_78__4, 
         camera_module_cache_ram_62__4, camera_module_cache_ram_46__4, 
         camera_module_cache_ram_30__4, camera_module_cache_ram_14__4, nx14740, 
         camera_module_cache_ram_253__4, camera_module_cache_ram_237__4, 
         camera_module_cache_ram_221__4, camera_module_cache_ram_205__4, 
         camera_module_cache_ram_189__4, camera_module_cache_ram_173__4, 
         camera_module_cache_ram_157__4, camera_module_cache_ram_141__4, nx14826, 
         camera_module_cache_ram_125__4, camera_module_cache_ram_109__4, 
         camera_module_cache_ram_93__4, camera_module_cache_ram_77__4, 
         camera_module_cache_ram_61__4, camera_module_cache_ram_45__4, 
         camera_module_cache_ram_29__4, camera_module_cache_ram_13__4, nx14904, 
         camera_module_cache_ram_252__4, camera_module_cache_ram_236__4, 
         camera_module_cache_ram_220__4, camera_module_cache_ram_204__4, 
         camera_module_cache_ram_188__4, camera_module_cache_ram_172__4, 
         camera_module_cache_ram_156__4, camera_module_cache_ram_140__4, nx14988, 
         camera_module_cache_ram_124__4, camera_module_cache_ram_108__4, 
         camera_module_cache_ram_92__4, camera_module_cache_ram_76__4, 
         camera_module_cache_ram_60__4, camera_module_cache_ram_44__4, 
         camera_module_cache_ram_28__4, camera_module_cache_ram_12__4, nx15066, 
         nx15076, camera_module_cache_ram_251__4, camera_module_cache_ram_235__4, 
         camera_module_cache_ram_219__4, camera_module_cache_ram_203__4, 
         camera_module_cache_ram_187__4, camera_module_cache_ram_171__4, 
         camera_module_cache_ram_155__4, camera_module_cache_ram_139__4, nx15154, 
         camera_module_cache_ram_123__4, camera_module_cache_ram_107__4, 
         camera_module_cache_ram_91__4, camera_module_cache_ram_75__4, 
         camera_module_cache_ram_59__4, camera_module_cache_ram_43__4, 
         camera_module_cache_ram_27__4, camera_module_cache_ram_11__4, nx15232, 
         camera_module_cache_ram_250__4, camera_module_cache_ram_234__4, 
         camera_module_cache_ram_218__4, camera_module_cache_ram_202__4, 
         camera_module_cache_ram_186__4, camera_module_cache_ram_170__4, 
         camera_module_cache_ram_154__4, camera_module_cache_ram_138__4, nx15316, 
         camera_module_cache_ram_122__4, camera_module_cache_ram_106__4, 
         camera_module_cache_ram_90__4, camera_module_cache_ram_74__4, 
         camera_module_cache_ram_58__4, camera_module_cache_ram_42__4, 
         camera_module_cache_ram_26__4, camera_module_cache_ram_10__4, nx15394, 
         camera_module_cache_ram_249__4, camera_module_cache_ram_233__4, 
         camera_module_cache_ram_217__4, camera_module_cache_ram_201__4, 
         camera_module_cache_ram_185__4, camera_module_cache_ram_169__4, 
         camera_module_cache_ram_153__4, camera_module_cache_ram_137__4, nx15480, 
         camera_module_cache_ram_121__4, camera_module_cache_ram_105__4, 
         camera_module_cache_ram_89__4, camera_module_cache_ram_73__4, 
         camera_module_cache_ram_57__4, camera_module_cache_ram_41__4, 
         camera_module_cache_ram_25__4, camera_module_cache_ram_9__4, nx15558, 
         camera_module_cache_ram_248__4, camera_module_cache_ram_232__4, 
         camera_module_cache_ram_216__4, camera_module_cache_ram_200__4, 
         camera_module_cache_ram_184__4, camera_module_cache_ram_168__4, 
         camera_module_cache_ram_152__4, camera_module_cache_ram_136__4, nx15642, 
         camera_module_cache_ram_120__4, camera_module_cache_ram_104__4, 
         camera_module_cache_ram_88__4, camera_module_cache_ram_72__4, 
         camera_module_cache_ram_56__4, camera_module_cache_ram_40__4, 
         camera_module_cache_ram_24__4, camera_module_cache_ram_8__4, nx15720, 
         nx15730, camera_module_cache_ram_247__4, camera_module_cache_ram_231__4, 
         camera_module_cache_ram_215__4, camera_module_cache_ram_199__4, 
         camera_module_cache_ram_183__4, camera_module_cache_ram_167__4, 
         camera_module_cache_ram_151__4, camera_module_cache_ram_135__4, nx15810, 
         camera_module_cache_ram_119__4, camera_module_cache_ram_103__4, 
         camera_module_cache_ram_87__4, camera_module_cache_ram_71__4, 
         camera_module_cache_ram_55__4, camera_module_cache_ram_39__4, 
         camera_module_cache_ram_23__4, camera_module_cache_ram_7__4, nx15888, 
         camera_module_cache_ram_246__4, camera_module_cache_ram_230__4, 
         camera_module_cache_ram_214__4, camera_module_cache_ram_198__4, 
         camera_module_cache_ram_182__4, camera_module_cache_ram_166__4, 
         camera_module_cache_ram_150__4, camera_module_cache_ram_134__4, nx15972, 
         camera_module_cache_ram_118__4, camera_module_cache_ram_102__4, 
         camera_module_cache_ram_86__4, camera_module_cache_ram_70__4, 
         camera_module_cache_ram_54__4, camera_module_cache_ram_38__4, 
         camera_module_cache_ram_22__4, camera_module_cache_ram_6__4, nx16050, 
         camera_module_cache_ram_245__4, camera_module_cache_ram_229__4, 
         camera_module_cache_ram_213__4, camera_module_cache_ram_197__4, 
         camera_module_cache_ram_181__4, camera_module_cache_ram_165__4, 
         camera_module_cache_ram_149__4, camera_module_cache_ram_133__4, nx16136, 
         camera_module_cache_ram_117__4, camera_module_cache_ram_101__4, 
         camera_module_cache_ram_85__4, camera_module_cache_ram_69__4, 
         camera_module_cache_ram_53__4, camera_module_cache_ram_37__4, 
         camera_module_cache_ram_21__4, camera_module_cache_ram_5__4, nx16214, 
         camera_module_cache_ram_244__4, camera_module_cache_ram_228__4, 
         camera_module_cache_ram_212__4, camera_module_cache_ram_196__4, 
         camera_module_cache_ram_180__4, camera_module_cache_ram_164__4, 
         camera_module_cache_ram_148__4, camera_module_cache_ram_132__4, nx16298, 
         camera_module_cache_ram_116__4, camera_module_cache_ram_100__4, 
         camera_module_cache_ram_84__4, camera_module_cache_ram_68__4, 
         camera_module_cache_ram_52__4, camera_module_cache_ram_36__4, 
         camera_module_cache_ram_20__4, camera_module_cache_ram_4__4, nx16376, 
         nx16386, camera_module_cache_ram_243__4, camera_module_cache_ram_227__4, 
         camera_module_cache_ram_211__4, camera_module_cache_ram_195__4, 
         camera_module_cache_ram_179__4, camera_module_cache_ram_163__4, 
         camera_module_cache_ram_147__4, camera_module_cache_ram_131__4, nx16464, 
         camera_module_cache_ram_115__4, camera_module_cache_ram_99__4, 
         camera_module_cache_ram_83__4, camera_module_cache_ram_67__4, 
         camera_module_cache_ram_51__4, camera_module_cache_ram_35__4, 
         camera_module_cache_ram_19__4, camera_module_cache_ram_3__4, nx16542, 
         camera_module_cache_ram_242__4, camera_module_cache_ram_226__4, 
         camera_module_cache_ram_210__4, camera_module_cache_ram_194__4, 
         camera_module_cache_ram_178__4, camera_module_cache_ram_162__4, 
         camera_module_cache_ram_146__4, camera_module_cache_ram_130__4, nx16626, 
         camera_module_cache_ram_114__4, camera_module_cache_ram_98__4, 
         camera_module_cache_ram_82__4, camera_module_cache_ram_66__4, 
         camera_module_cache_ram_50__4, camera_module_cache_ram_34__4, 
         camera_module_cache_ram_18__4, camera_module_cache_ram_2__4, nx16704, 
         camera_module_cache_ram_241__4, camera_module_cache_ram_225__4, 
         camera_module_cache_ram_209__4, camera_module_cache_ram_193__4, 
         camera_module_cache_ram_177__4, camera_module_cache_ram_161__4, 
         camera_module_cache_ram_145__4, camera_module_cache_ram_129__4, nx16790, 
         camera_module_cache_ram_113__4, camera_module_cache_ram_97__4, 
         camera_module_cache_ram_81__4, camera_module_cache_ram_65__4, 
         camera_module_cache_ram_49__4, camera_module_cache_ram_33__4, 
         camera_module_cache_ram_17__4, camera_module_cache_ram_1__4, nx16868, 
         camera_module_cache_ram_240__4, camera_module_cache_ram_224__4, 
         camera_module_cache_ram_208__4, camera_module_cache_ram_192__4, 
         camera_module_cache_ram_176__4, camera_module_cache_ram_160__4, 
         camera_module_cache_ram_144__4, camera_module_cache_ram_128__4, nx16952, 
         camera_module_cache_ram_112__4, camera_module_cache_ram_96__4, 
         camera_module_cache_ram_80__4, camera_module_cache_ram_64__4, 
         camera_module_cache_ram_48__4, camera_module_cache_ram_32__4, 
         camera_module_cache_ram_16__4, camera_module_cache_ram_0__4, nx17030, 
         nx17040, nx17060, nx17068, camera_module_algo_module_pixel_value_5, 
         camera_module_cache_ram_255__5, nx17098, nx17108, nx17120, nx17124, 
         nx17130, nx17140, nx17152, nx17156, nx17168, nx17180, nx17184, nx17196, 
         camera_module_cache_ram_239__5, camera_module_cache_ram_223__5, 
         camera_module_cache_ram_207__5, camera_module_cache_ram_191__5, 
         camera_module_cache_ram_175__5, camera_module_cache_ram_159__5, 
         camera_module_cache_ram_143__5, nx17274, camera_module_cache_ram_127__5, 
         camera_module_cache_ram_111__5, camera_module_cache_ram_95__5, 
         camera_module_cache_ram_79__5, camera_module_cache_ram_63__5, 
         camera_module_cache_ram_47__5, camera_module_cache_ram_31__5, 
         camera_module_cache_ram_15__5, nx17352, camera_module_cache_ram_254__5, 
         camera_module_cache_ram_238__5, camera_module_cache_ram_222__5, 
         camera_module_cache_ram_206__5, camera_module_cache_ram_190__5, 
         camera_module_cache_ram_174__5, camera_module_cache_ram_158__5, 
         camera_module_cache_ram_142__5, nx17436, camera_module_cache_ram_126__5, 
         camera_module_cache_ram_110__5, camera_module_cache_ram_94__5, 
         camera_module_cache_ram_78__5, camera_module_cache_ram_62__5, 
         camera_module_cache_ram_46__5, camera_module_cache_ram_30__5, 
         camera_module_cache_ram_14__5, nx17514, camera_module_cache_ram_253__5, 
         camera_module_cache_ram_237__5, camera_module_cache_ram_221__5, 
         camera_module_cache_ram_205__5, camera_module_cache_ram_189__5, 
         camera_module_cache_ram_173__5, camera_module_cache_ram_157__5, 
         camera_module_cache_ram_141__5, nx17600, camera_module_cache_ram_125__5, 
         camera_module_cache_ram_109__5, camera_module_cache_ram_93__5, 
         camera_module_cache_ram_77__5, camera_module_cache_ram_61__5, 
         camera_module_cache_ram_45__5, camera_module_cache_ram_29__5, 
         camera_module_cache_ram_13__5, nx17678, camera_module_cache_ram_252__5, 
         camera_module_cache_ram_236__5, camera_module_cache_ram_220__5, 
         camera_module_cache_ram_204__5, camera_module_cache_ram_188__5, 
         camera_module_cache_ram_172__5, camera_module_cache_ram_156__5, 
         camera_module_cache_ram_140__5, nx17762, camera_module_cache_ram_124__5, 
         camera_module_cache_ram_108__5, camera_module_cache_ram_92__5, 
         camera_module_cache_ram_76__5, camera_module_cache_ram_60__5, 
         camera_module_cache_ram_44__5, camera_module_cache_ram_28__5, 
         camera_module_cache_ram_12__5, nx17840, nx17850, 
         camera_module_cache_ram_251__5, camera_module_cache_ram_235__5, 
         camera_module_cache_ram_219__5, camera_module_cache_ram_203__5, 
         camera_module_cache_ram_187__5, camera_module_cache_ram_171__5, 
         camera_module_cache_ram_155__5, camera_module_cache_ram_139__5, nx17928, 
         camera_module_cache_ram_123__5, camera_module_cache_ram_107__5, 
         camera_module_cache_ram_91__5, camera_module_cache_ram_75__5, 
         camera_module_cache_ram_59__5, camera_module_cache_ram_43__5, 
         camera_module_cache_ram_27__5, camera_module_cache_ram_11__5, nx18006, 
         camera_module_cache_ram_250__5, camera_module_cache_ram_234__5, 
         camera_module_cache_ram_218__5, camera_module_cache_ram_202__5, 
         camera_module_cache_ram_186__5, camera_module_cache_ram_170__5, 
         camera_module_cache_ram_154__5, camera_module_cache_ram_138__5, nx18090, 
         camera_module_cache_ram_122__5, camera_module_cache_ram_106__5, 
         camera_module_cache_ram_90__5, camera_module_cache_ram_74__5, 
         camera_module_cache_ram_58__5, camera_module_cache_ram_42__5, 
         camera_module_cache_ram_26__5, camera_module_cache_ram_10__5, nx18168, 
         camera_module_cache_ram_249__5, camera_module_cache_ram_233__5, 
         camera_module_cache_ram_217__5, camera_module_cache_ram_201__5, 
         camera_module_cache_ram_185__5, camera_module_cache_ram_169__5, 
         camera_module_cache_ram_153__5, camera_module_cache_ram_137__5, nx18254, 
         camera_module_cache_ram_121__5, camera_module_cache_ram_105__5, 
         camera_module_cache_ram_89__5, camera_module_cache_ram_73__5, 
         camera_module_cache_ram_57__5, camera_module_cache_ram_41__5, 
         camera_module_cache_ram_25__5, camera_module_cache_ram_9__5, nx18332, 
         camera_module_cache_ram_248__5, camera_module_cache_ram_232__5, 
         camera_module_cache_ram_216__5, camera_module_cache_ram_200__5, 
         camera_module_cache_ram_184__5, camera_module_cache_ram_168__5, 
         camera_module_cache_ram_152__5, camera_module_cache_ram_136__5, nx18416, 
         camera_module_cache_ram_120__5, camera_module_cache_ram_104__5, 
         camera_module_cache_ram_88__5, camera_module_cache_ram_72__5, 
         camera_module_cache_ram_56__5, camera_module_cache_ram_40__5, 
         camera_module_cache_ram_24__5, camera_module_cache_ram_8__5, nx18494, 
         nx18504, camera_module_cache_ram_247__5, camera_module_cache_ram_231__5, 
         camera_module_cache_ram_215__5, camera_module_cache_ram_199__5, 
         camera_module_cache_ram_183__5, camera_module_cache_ram_167__5, 
         camera_module_cache_ram_151__5, camera_module_cache_ram_135__5, nx18584, 
         camera_module_cache_ram_119__5, camera_module_cache_ram_103__5, 
         camera_module_cache_ram_87__5, camera_module_cache_ram_71__5, 
         camera_module_cache_ram_55__5, camera_module_cache_ram_39__5, 
         camera_module_cache_ram_23__5, camera_module_cache_ram_7__5, nx18662, 
         camera_module_cache_ram_246__5, camera_module_cache_ram_230__5, 
         camera_module_cache_ram_214__5, camera_module_cache_ram_198__5, 
         camera_module_cache_ram_182__5, camera_module_cache_ram_166__5, 
         camera_module_cache_ram_150__5, camera_module_cache_ram_134__5, nx18746, 
         camera_module_cache_ram_118__5, camera_module_cache_ram_102__5, 
         camera_module_cache_ram_86__5, camera_module_cache_ram_70__5, 
         camera_module_cache_ram_54__5, camera_module_cache_ram_38__5, 
         camera_module_cache_ram_22__5, camera_module_cache_ram_6__5, nx18824, 
         camera_module_cache_ram_245__5, camera_module_cache_ram_229__5, 
         camera_module_cache_ram_213__5, camera_module_cache_ram_197__5, 
         camera_module_cache_ram_181__5, camera_module_cache_ram_165__5, 
         camera_module_cache_ram_149__5, camera_module_cache_ram_133__5, nx18910, 
         camera_module_cache_ram_117__5, camera_module_cache_ram_101__5, 
         camera_module_cache_ram_85__5, camera_module_cache_ram_69__5, 
         camera_module_cache_ram_53__5, camera_module_cache_ram_37__5, 
         camera_module_cache_ram_21__5, camera_module_cache_ram_5__5, nx18988, 
         camera_module_cache_ram_244__5, camera_module_cache_ram_228__5, 
         camera_module_cache_ram_212__5, camera_module_cache_ram_196__5, 
         camera_module_cache_ram_180__5, camera_module_cache_ram_164__5, 
         camera_module_cache_ram_148__5, camera_module_cache_ram_132__5, nx19072, 
         camera_module_cache_ram_116__5, camera_module_cache_ram_100__5, 
         camera_module_cache_ram_84__5, camera_module_cache_ram_68__5, 
         camera_module_cache_ram_52__5, camera_module_cache_ram_36__5, 
         camera_module_cache_ram_20__5, camera_module_cache_ram_4__5, nx19150, 
         nx19160, camera_module_cache_ram_243__5, camera_module_cache_ram_227__5, 
         camera_module_cache_ram_211__5, camera_module_cache_ram_195__5, 
         camera_module_cache_ram_179__5, camera_module_cache_ram_163__5, 
         camera_module_cache_ram_147__5, camera_module_cache_ram_131__5, nx19238, 
         camera_module_cache_ram_115__5, camera_module_cache_ram_99__5, 
         camera_module_cache_ram_83__5, camera_module_cache_ram_67__5, 
         camera_module_cache_ram_51__5, camera_module_cache_ram_35__5, 
         camera_module_cache_ram_19__5, camera_module_cache_ram_3__5, nx19316, 
         camera_module_cache_ram_242__5, camera_module_cache_ram_226__5, 
         camera_module_cache_ram_210__5, camera_module_cache_ram_194__5, 
         camera_module_cache_ram_178__5, camera_module_cache_ram_162__5, 
         camera_module_cache_ram_146__5, camera_module_cache_ram_130__5, nx19400, 
         camera_module_cache_ram_114__5, camera_module_cache_ram_98__5, 
         camera_module_cache_ram_82__5, camera_module_cache_ram_66__5, 
         camera_module_cache_ram_50__5, camera_module_cache_ram_34__5, 
         camera_module_cache_ram_18__5, camera_module_cache_ram_2__5, nx19478, 
         camera_module_cache_ram_241__5, camera_module_cache_ram_225__5, 
         camera_module_cache_ram_209__5, camera_module_cache_ram_193__5, 
         camera_module_cache_ram_177__5, camera_module_cache_ram_161__5, 
         camera_module_cache_ram_145__5, camera_module_cache_ram_129__5, nx19564, 
         camera_module_cache_ram_113__5, camera_module_cache_ram_97__5, 
         camera_module_cache_ram_81__5, camera_module_cache_ram_65__5, 
         camera_module_cache_ram_49__5, camera_module_cache_ram_33__5, 
         camera_module_cache_ram_17__5, camera_module_cache_ram_1__5, nx19642, 
         camera_module_cache_ram_240__5, camera_module_cache_ram_224__5, 
         camera_module_cache_ram_208__5, camera_module_cache_ram_192__5, 
         camera_module_cache_ram_176__5, camera_module_cache_ram_160__5, 
         camera_module_cache_ram_144__5, camera_module_cache_ram_128__5, nx19726, 
         camera_module_cache_ram_112__5, camera_module_cache_ram_96__5, 
         camera_module_cache_ram_80__5, camera_module_cache_ram_64__5, 
         camera_module_cache_ram_48__5, camera_module_cache_ram_32__5, 
         camera_module_cache_ram_16__5, camera_module_cache_ram_0__5, nx19804, 
         nx19814, nx19826, nx19834, nx19850, 
         camera_module_algo_module_pixel_value_6, camera_module_cache_ram_255__6, 
         nx19872, nx19882, nx19894, nx19898, nx19904, nx19914, nx19926, nx19930, 
         nx19942, nx19954, nx19958, nx19970, camera_module_cache_ram_239__6, 
         camera_module_cache_ram_223__6, camera_module_cache_ram_207__6, 
         camera_module_cache_ram_191__6, camera_module_cache_ram_175__6, 
         camera_module_cache_ram_159__6, camera_module_cache_ram_143__6, nx20048, 
         camera_module_cache_ram_127__6, camera_module_cache_ram_111__6, 
         camera_module_cache_ram_95__6, camera_module_cache_ram_79__6, 
         camera_module_cache_ram_63__6, camera_module_cache_ram_47__6, 
         camera_module_cache_ram_31__6, camera_module_cache_ram_15__6, nx20126, 
         camera_module_cache_ram_254__6, camera_module_cache_ram_238__6, 
         camera_module_cache_ram_222__6, camera_module_cache_ram_206__6, 
         camera_module_cache_ram_190__6, camera_module_cache_ram_174__6, 
         camera_module_cache_ram_158__6, camera_module_cache_ram_142__6, nx20210, 
         camera_module_cache_ram_126__6, camera_module_cache_ram_110__6, 
         camera_module_cache_ram_94__6, camera_module_cache_ram_78__6, 
         camera_module_cache_ram_62__6, camera_module_cache_ram_46__6, 
         camera_module_cache_ram_30__6, camera_module_cache_ram_14__6, nx20288, 
         camera_module_cache_ram_253__6, camera_module_cache_ram_237__6, 
         camera_module_cache_ram_221__6, camera_module_cache_ram_205__6, 
         camera_module_cache_ram_189__6, camera_module_cache_ram_173__6, 
         camera_module_cache_ram_157__6, camera_module_cache_ram_141__6, nx20374, 
         camera_module_cache_ram_125__6, camera_module_cache_ram_109__6, 
         camera_module_cache_ram_93__6, camera_module_cache_ram_77__6, 
         camera_module_cache_ram_61__6, camera_module_cache_ram_45__6, 
         camera_module_cache_ram_29__6, camera_module_cache_ram_13__6, nx20452, 
         camera_module_cache_ram_252__6, camera_module_cache_ram_236__6, 
         camera_module_cache_ram_220__6, camera_module_cache_ram_204__6, 
         camera_module_cache_ram_188__6, camera_module_cache_ram_172__6, 
         camera_module_cache_ram_156__6, camera_module_cache_ram_140__6, nx20536, 
         camera_module_cache_ram_124__6, camera_module_cache_ram_108__6, 
         camera_module_cache_ram_92__6, camera_module_cache_ram_76__6, 
         camera_module_cache_ram_60__6, camera_module_cache_ram_44__6, 
         camera_module_cache_ram_28__6, camera_module_cache_ram_12__6, nx20614, 
         nx20624, camera_module_cache_ram_251__6, camera_module_cache_ram_235__6, 
         camera_module_cache_ram_219__6, camera_module_cache_ram_203__6, 
         camera_module_cache_ram_187__6, camera_module_cache_ram_171__6, 
         camera_module_cache_ram_155__6, camera_module_cache_ram_139__6, nx20702, 
         camera_module_cache_ram_123__6, camera_module_cache_ram_107__6, 
         camera_module_cache_ram_91__6, camera_module_cache_ram_75__6, 
         camera_module_cache_ram_59__6, camera_module_cache_ram_43__6, 
         camera_module_cache_ram_27__6, camera_module_cache_ram_11__6, nx20780, 
         camera_module_cache_ram_250__6, camera_module_cache_ram_234__6, 
         camera_module_cache_ram_218__6, camera_module_cache_ram_202__6, 
         camera_module_cache_ram_186__6, camera_module_cache_ram_170__6, 
         camera_module_cache_ram_154__6, camera_module_cache_ram_138__6, nx20864, 
         camera_module_cache_ram_122__6, camera_module_cache_ram_106__6, 
         camera_module_cache_ram_90__6, camera_module_cache_ram_74__6, 
         camera_module_cache_ram_58__6, camera_module_cache_ram_42__6, 
         camera_module_cache_ram_26__6, camera_module_cache_ram_10__6, nx20942, 
         camera_module_cache_ram_249__6, camera_module_cache_ram_233__6, 
         camera_module_cache_ram_217__6, camera_module_cache_ram_201__6, 
         camera_module_cache_ram_185__6, camera_module_cache_ram_169__6, 
         camera_module_cache_ram_153__6, camera_module_cache_ram_137__6, nx21028, 
         camera_module_cache_ram_121__6, camera_module_cache_ram_105__6, 
         camera_module_cache_ram_89__6, camera_module_cache_ram_73__6, 
         camera_module_cache_ram_57__6, camera_module_cache_ram_41__6, 
         camera_module_cache_ram_25__6, camera_module_cache_ram_9__6, nx21106, 
         camera_module_cache_ram_248__6, camera_module_cache_ram_232__6, 
         camera_module_cache_ram_216__6, camera_module_cache_ram_200__6, 
         camera_module_cache_ram_184__6, camera_module_cache_ram_168__6, 
         camera_module_cache_ram_152__6, camera_module_cache_ram_136__6, nx21190, 
         camera_module_cache_ram_120__6, camera_module_cache_ram_104__6, 
         camera_module_cache_ram_88__6, camera_module_cache_ram_72__6, 
         camera_module_cache_ram_56__6, camera_module_cache_ram_40__6, 
         camera_module_cache_ram_24__6, camera_module_cache_ram_8__6, nx21268, 
         nx21278, camera_module_cache_ram_247__6, camera_module_cache_ram_231__6, 
         camera_module_cache_ram_215__6, camera_module_cache_ram_199__6, 
         camera_module_cache_ram_183__6, camera_module_cache_ram_167__6, 
         camera_module_cache_ram_151__6, camera_module_cache_ram_135__6, nx21358, 
         camera_module_cache_ram_119__6, camera_module_cache_ram_103__6, 
         camera_module_cache_ram_87__6, camera_module_cache_ram_71__6, 
         camera_module_cache_ram_55__6, camera_module_cache_ram_39__6, 
         camera_module_cache_ram_23__6, camera_module_cache_ram_7__6, nx21436, 
         camera_module_cache_ram_246__6, camera_module_cache_ram_230__6, 
         camera_module_cache_ram_214__6, camera_module_cache_ram_198__6, 
         camera_module_cache_ram_182__6, camera_module_cache_ram_166__6, 
         camera_module_cache_ram_150__6, camera_module_cache_ram_134__6, nx21520, 
         camera_module_cache_ram_118__6, camera_module_cache_ram_102__6, 
         camera_module_cache_ram_86__6, camera_module_cache_ram_70__6, 
         camera_module_cache_ram_54__6, camera_module_cache_ram_38__6, 
         camera_module_cache_ram_22__6, camera_module_cache_ram_6__6, nx21598, 
         camera_module_cache_ram_245__6, camera_module_cache_ram_229__6, 
         camera_module_cache_ram_213__6, camera_module_cache_ram_197__6, 
         camera_module_cache_ram_181__6, camera_module_cache_ram_165__6, 
         camera_module_cache_ram_149__6, camera_module_cache_ram_133__6, nx21684, 
         camera_module_cache_ram_117__6, camera_module_cache_ram_101__6, 
         camera_module_cache_ram_85__6, camera_module_cache_ram_69__6, 
         camera_module_cache_ram_53__6, camera_module_cache_ram_37__6, 
         camera_module_cache_ram_21__6, camera_module_cache_ram_5__6, nx21762, 
         camera_module_cache_ram_244__6, camera_module_cache_ram_228__6, 
         camera_module_cache_ram_212__6, camera_module_cache_ram_196__6, 
         camera_module_cache_ram_180__6, camera_module_cache_ram_164__6, 
         camera_module_cache_ram_148__6, camera_module_cache_ram_132__6, nx21846, 
         camera_module_cache_ram_116__6, camera_module_cache_ram_100__6, 
         camera_module_cache_ram_84__6, camera_module_cache_ram_68__6, 
         camera_module_cache_ram_52__6, camera_module_cache_ram_36__6, 
         camera_module_cache_ram_20__6, camera_module_cache_ram_4__6, nx21924, 
         nx21934, camera_module_cache_ram_243__6, camera_module_cache_ram_227__6, 
         camera_module_cache_ram_211__6, camera_module_cache_ram_195__6, 
         camera_module_cache_ram_179__6, camera_module_cache_ram_163__6, 
         camera_module_cache_ram_147__6, camera_module_cache_ram_131__6, nx22012, 
         camera_module_cache_ram_115__6, camera_module_cache_ram_99__6, 
         camera_module_cache_ram_83__6, camera_module_cache_ram_67__6, 
         camera_module_cache_ram_51__6, camera_module_cache_ram_35__6, 
         camera_module_cache_ram_19__6, camera_module_cache_ram_3__6, nx22090, 
         camera_module_cache_ram_242__6, camera_module_cache_ram_226__6, 
         camera_module_cache_ram_210__6, camera_module_cache_ram_194__6, 
         camera_module_cache_ram_178__6, camera_module_cache_ram_162__6, 
         camera_module_cache_ram_146__6, camera_module_cache_ram_130__6, nx22174, 
         camera_module_cache_ram_114__6, camera_module_cache_ram_98__6, 
         camera_module_cache_ram_82__6, camera_module_cache_ram_66__6, 
         camera_module_cache_ram_50__6, camera_module_cache_ram_34__6, 
         camera_module_cache_ram_18__6, camera_module_cache_ram_2__6, nx22252, 
         camera_module_cache_ram_241__6, camera_module_cache_ram_225__6, 
         camera_module_cache_ram_209__6, camera_module_cache_ram_193__6, 
         camera_module_cache_ram_177__6, camera_module_cache_ram_161__6, 
         camera_module_cache_ram_145__6, camera_module_cache_ram_129__6, nx22338, 
         camera_module_cache_ram_113__6, camera_module_cache_ram_97__6, 
         camera_module_cache_ram_81__6, camera_module_cache_ram_65__6, 
         camera_module_cache_ram_49__6, camera_module_cache_ram_33__6, 
         camera_module_cache_ram_17__6, camera_module_cache_ram_1__6, nx22416, 
         camera_module_cache_ram_240__6, camera_module_cache_ram_224__6, 
         camera_module_cache_ram_208__6, camera_module_cache_ram_192__6, 
         camera_module_cache_ram_176__6, camera_module_cache_ram_160__6, 
         camera_module_cache_ram_144__6, camera_module_cache_ram_128__6, nx22500, 
         camera_module_cache_ram_112__6, camera_module_cache_ram_96__6, 
         camera_module_cache_ram_80__6, camera_module_cache_ram_64__6, 
         camera_module_cache_ram_48__6, camera_module_cache_ram_32__6, 
         camera_module_cache_ram_16__6, camera_module_cache_ram_0__6, nx22578, 
         nx22588, nx22608, nx22616, camera_module_algo_module_pixel_value_7, 
         camera_module_cache_ram_255__7, nx22646, nx22656, nx22668, nx22672, 
         nx22678, nx22688, nx22700, nx22704, nx22716, nx22728, nx22732, nx22744, 
         camera_module_cache_ram_239__7, camera_module_cache_ram_223__7, 
         camera_module_cache_ram_207__7, camera_module_cache_ram_191__7, 
         camera_module_cache_ram_175__7, camera_module_cache_ram_159__7, 
         camera_module_cache_ram_143__7, nx22822, camera_module_cache_ram_127__7, 
         camera_module_cache_ram_111__7, camera_module_cache_ram_95__7, 
         camera_module_cache_ram_79__7, camera_module_cache_ram_63__7, 
         camera_module_cache_ram_47__7, camera_module_cache_ram_31__7, 
         camera_module_cache_ram_15__7, nx22900, camera_module_cache_ram_254__7, 
         camera_module_cache_ram_238__7, camera_module_cache_ram_222__7, 
         camera_module_cache_ram_206__7, camera_module_cache_ram_190__7, 
         camera_module_cache_ram_174__7, camera_module_cache_ram_158__7, 
         camera_module_cache_ram_142__7, nx22984, camera_module_cache_ram_126__7, 
         camera_module_cache_ram_110__7, camera_module_cache_ram_94__7, 
         camera_module_cache_ram_78__7, camera_module_cache_ram_62__7, 
         camera_module_cache_ram_46__7, camera_module_cache_ram_30__7, 
         camera_module_cache_ram_14__7, nx23062, camera_module_cache_ram_253__7, 
         camera_module_cache_ram_237__7, camera_module_cache_ram_221__7, 
         camera_module_cache_ram_205__7, camera_module_cache_ram_189__7, 
         camera_module_cache_ram_173__7, camera_module_cache_ram_157__7, 
         camera_module_cache_ram_141__7, nx23148, camera_module_cache_ram_125__7, 
         camera_module_cache_ram_109__7, camera_module_cache_ram_93__7, 
         camera_module_cache_ram_77__7, camera_module_cache_ram_61__7, 
         camera_module_cache_ram_45__7, camera_module_cache_ram_29__7, 
         camera_module_cache_ram_13__7, nx23226, camera_module_cache_ram_252__7, 
         camera_module_cache_ram_236__7, camera_module_cache_ram_220__7, 
         camera_module_cache_ram_204__7, camera_module_cache_ram_188__7, 
         camera_module_cache_ram_172__7, camera_module_cache_ram_156__7, 
         camera_module_cache_ram_140__7, nx23310, camera_module_cache_ram_124__7, 
         camera_module_cache_ram_108__7, camera_module_cache_ram_92__7, 
         camera_module_cache_ram_76__7, camera_module_cache_ram_60__7, 
         camera_module_cache_ram_44__7, camera_module_cache_ram_28__7, 
         camera_module_cache_ram_12__7, nx23388, nx23398, 
         camera_module_cache_ram_251__7, camera_module_cache_ram_235__7, 
         camera_module_cache_ram_219__7, camera_module_cache_ram_203__7, 
         camera_module_cache_ram_187__7, camera_module_cache_ram_171__7, 
         camera_module_cache_ram_155__7, camera_module_cache_ram_139__7, nx23476, 
         camera_module_cache_ram_123__7, camera_module_cache_ram_107__7, 
         camera_module_cache_ram_91__7, camera_module_cache_ram_75__7, 
         camera_module_cache_ram_59__7, camera_module_cache_ram_43__7, 
         camera_module_cache_ram_27__7, camera_module_cache_ram_11__7, nx23554, 
         camera_module_cache_ram_250__7, camera_module_cache_ram_234__7, 
         camera_module_cache_ram_218__7, camera_module_cache_ram_202__7, 
         camera_module_cache_ram_186__7, camera_module_cache_ram_170__7, 
         camera_module_cache_ram_154__7, camera_module_cache_ram_138__7, nx23638, 
         camera_module_cache_ram_122__7, camera_module_cache_ram_106__7, 
         camera_module_cache_ram_90__7, camera_module_cache_ram_74__7, 
         camera_module_cache_ram_58__7, camera_module_cache_ram_42__7, 
         camera_module_cache_ram_26__7, camera_module_cache_ram_10__7, nx23716, 
         camera_module_cache_ram_249__7, camera_module_cache_ram_233__7, 
         camera_module_cache_ram_217__7, camera_module_cache_ram_201__7, 
         camera_module_cache_ram_185__7, camera_module_cache_ram_169__7, 
         camera_module_cache_ram_153__7, camera_module_cache_ram_137__7, nx23802, 
         camera_module_cache_ram_121__7, camera_module_cache_ram_105__7, 
         camera_module_cache_ram_89__7, camera_module_cache_ram_73__7, 
         camera_module_cache_ram_57__7, camera_module_cache_ram_41__7, 
         camera_module_cache_ram_25__7, camera_module_cache_ram_9__7, nx23880, 
         camera_module_cache_ram_248__7, camera_module_cache_ram_232__7, 
         camera_module_cache_ram_216__7, camera_module_cache_ram_200__7, 
         camera_module_cache_ram_184__7, camera_module_cache_ram_168__7, 
         camera_module_cache_ram_152__7, camera_module_cache_ram_136__7, nx23964, 
         camera_module_cache_ram_120__7, camera_module_cache_ram_104__7, 
         camera_module_cache_ram_88__7, camera_module_cache_ram_72__7, 
         camera_module_cache_ram_56__7, camera_module_cache_ram_40__7, 
         camera_module_cache_ram_24__7, camera_module_cache_ram_8__7, nx24042, 
         nx24052, camera_module_cache_ram_247__7, camera_module_cache_ram_231__7, 
         camera_module_cache_ram_215__7, camera_module_cache_ram_199__7, 
         camera_module_cache_ram_183__7, camera_module_cache_ram_167__7, 
         camera_module_cache_ram_151__7, camera_module_cache_ram_135__7, nx24132, 
         camera_module_cache_ram_119__7, camera_module_cache_ram_103__7, 
         camera_module_cache_ram_87__7, camera_module_cache_ram_71__7, 
         camera_module_cache_ram_55__7, camera_module_cache_ram_39__7, 
         camera_module_cache_ram_23__7, camera_module_cache_ram_7__7, nx24210, 
         camera_module_cache_ram_246__7, camera_module_cache_ram_230__7, 
         camera_module_cache_ram_214__7, camera_module_cache_ram_198__7, 
         camera_module_cache_ram_182__7, camera_module_cache_ram_166__7, 
         camera_module_cache_ram_150__7, camera_module_cache_ram_134__7, nx24294, 
         camera_module_cache_ram_118__7, camera_module_cache_ram_102__7, 
         camera_module_cache_ram_86__7, camera_module_cache_ram_70__7, 
         camera_module_cache_ram_54__7, camera_module_cache_ram_38__7, 
         camera_module_cache_ram_22__7, camera_module_cache_ram_6__7, nx24372, 
         camera_module_cache_ram_245__7, camera_module_cache_ram_229__7, 
         camera_module_cache_ram_213__7, camera_module_cache_ram_197__7, 
         camera_module_cache_ram_181__7, camera_module_cache_ram_165__7, 
         camera_module_cache_ram_149__7, camera_module_cache_ram_133__7, nx24458, 
         camera_module_cache_ram_117__7, camera_module_cache_ram_101__7, 
         camera_module_cache_ram_85__7, camera_module_cache_ram_69__7, 
         camera_module_cache_ram_53__7, camera_module_cache_ram_37__7, 
         camera_module_cache_ram_21__7, camera_module_cache_ram_5__7, nx24536, 
         camera_module_cache_ram_244__7, camera_module_cache_ram_228__7, 
         camera_module_cache_ram_212__7, camera_module_cache_ram_196__7, 
         camera_module_cache_ram_180__7, camera_module_cache_ram_164__7, 
         camera_module_cache_ram_148__7, camera_module_cache_ram_132__7, nx24620, 
         camera_module_cache_ram_116__7, camera_module_cache_ram_100__7, 
         camera_module_cache_ram_84__7, camera_module_cache_ram_68__7, 
         camera_module_cache_ram_52__7, camera_module_cache_ram_36__7, 
         camera_module_cache_ram_20__7, camera_module_cache_ram_4__7, nx24698, 
         nx24708, camera_module_cache_ram_243__7, camera_module_cache_ram_227__7, 
         camera_module_cache_ram_211__7, camera_module_cache_ram_195__7, 
         camera_module_cache_ram_179__7, camera_module_cache_ram_163__7, 
         camera_module_cache_ram_147__7, camera_module_cache_ram_131__7, nx24786, 
         camera_module_cache_ram_115__7, camera_module_cache_ram_99__7, 
         camera_module_cache_ram_83__7, camera_module_cache_ram_67__7, 
         camera_module_cache_ram_51__7, camera_module_cache_ram_35__7, 
         camera_module_cache_ram_19__7, camera_module_cache_ram_3__7, nx24864, 
         camera_module_cache_ram_242__7, camera_module_cache_ram_226__7, 
         camera_module_cache_ram_210__7, camera_module_cache_ram_194__7, 
         camera_module_cache_ram_178__7, camera_module_cache_ram_162__7, 
         camera_module_cache_ram_146__7, camera_module_cache_ram_130__7, nx24948, 
         camera_module_cache_ram_114__7, camera_module_cache_ram_98__7, 
         camera_module_cache_ram_82__7, camera_module_cache_ram_66__7, 
         camera_module_cache_ram_50__7, camera_module_cache_ram_34__7, 
         camera_module_cache_ram_18__7, camera_module_cache_ram_2__7, nx25026, 
         camera_module_cache_ram_241__7, camera_module_cache_ram_225__7, 
         camera_module_cache_ram_209__7, camera_module_cache_ram_193__7, 
         camera_module_cache_ram_177__7, camera_module_cache_ram_161__7, 
         camera_module_cache_ram_145__7, camera_module_cache_ram_129__7, nx25112, 
         camera_module_cache_ram_113__7, camera_module_cache_ram_97__7, 
         camera_module_cache_ram_81__7, camera_module_cache_ram_65__7, 
         camera_module_cache_ram_49__7, camera_module_cache_ram_33__7, 
         camera_module_cache_ram_17__7, camera_module_cache_ram_1__7, nx25190, 
         camera_module_cache_ram_240__7, camera_module_cache_ram_224__7, 
         camera_module_cache_ram_208__7, camera_module_cache_ram_192__7, 
         camera_module_cache_ram_176__7, camera_module_cache_ram_160__7, 
         camera_module_cache_ram_144__7, camera_module_cache_ram_128__7, nx25274, 
         camera_module_cache_ram_112__7, camera_module_cache_ram_96__7, 
         camera_module_cache_ram_80__7, camera_module_cache_ram_64__7, 
         camera_module_cache_ram_48__7, camera_module_cache_ram_32__7, 
         camera_module_cache_ram_16__7, camera_module_cache_ram_0__7, nx25352, 
         nx25362, nx25374, nx25382, nx25398, nx25406, nx25414, nx25422, nx25432, 
         nx25434, nx25436, nx25438, nx25446, nx25454, nx25468, 
         camera_module_algo_module_current_cont_value_1, 
         camera_module_algo_module_Addout_value_1, nx910, nx25470, nx25478, 
         nx25492, camera_module_algo_module_diff_value_1, nx25508, nx25520, 
         nx25528, camera_module_algo_module_current_cont_value_2, 
         camera_module_algo_module_Addout_value_2, nx25552, nx25566, 
         camera_module_algo_module_diff_value_2, nx25580, nx25582, nx25584, 
         nx25586, nx25594, nx25602, nx25616, 
         camera_module_algo_module_current_cont_value_3, 
         camera_module_algo_module_Addout_value_3, nx913, nx25618, nx25626, 
         nx25640, camera_module_algo_module_diff_value_3, nx25656, nx25668, 
         nx25676, camera_module_algo_module_current_cont_value_4, 
         camera_module_algo_module_Addout_value_4, nx25700, nx25714, 
         camera_module_algo_module_diff_value_4, nx25728, nx25730, nx25732, 
         nx25734, nx25742, nx25750, nx25764, 
         camera_module_algo_module_current_cont_value_5, 
         camera_module_algo_module_Addout_value_5, nx917, nx25766, nx25774, 
         nx25788, camera_module_algo_module_diff_value_5, nx25804, nx25816, 
         nx25824, camera_module_algo_module_current_cont_value_6, 
         camera_module_algo_module_Addout_value_6, nx25848, nx25862, 
         camera_module_algo_module_diff_value_6, nx25876, nx25878, nx25880, 
         nx25882, nx25890, nx25898, nx25912, 
         camera_module_algo_module_current_cont_value_7, 
         camera_module_algo_module_Addout_value_7, nx921, nx25914, nx25922, 
         nx25936, camera_module_algo_module_diff_value_7, nx25952, nx25964, 
         nx25972, camera_module_algo_module_current_cont_value_8, 
         camera_module_algo_module_Addout_value_8, nx25996, nx26010, 
         camera_module_algo_module_diff_value_8, nx26024, nx26026, nx26028, 
         nx26030, nx26038, nx26046, nx26060, 
         camera_module_algo_module_current_cont_value_9, 
         camera_module_algo_module_Addout_value_9, nx925, nx26062, nx26070, 
         nx26084, camera_module_algo_module_diff_value_9, nx26100, nx26116, 
         camera_module_algo_module_current_cont_value_10, 
         camera_module_algo_module_Addout_value_10, nx26144, nx26158, nx26172, 
         nx26174, nx26176, nx26190, nx26208, 
         camera_module_algo_module_current_cont_value_11, 
         camera_module_algo_module_Addout_value_11, nx929, nx26210, nx26218, 
         nx26232, camera_module_algo_module_diff_value_11, nx26248, nx26264, 
         camera_module_algo_module_current_cont_value_12, 
         camera_module_algo_module_Addout_value_12, nx26292, nx26306, nx26320, 
         nx26322, nx26324, nx26338, nx26356, 
         camera_module_algo_module_current_cont_value_13, 
         camera_module_algo_module_Addout_value_13, nx933, nx26358, nx26366, 
         nx26380, camera_module_algo_module_diff_value_13, nx26396, nx26412, 
         camera_module_algo_module_current_cont_value_14, 
         camera_module_algo_module_Addout_value_14, nx26440, nx26454, nx26468, 
         nx26470, nx26472, nx26486, nx26504, 
         camera_module_algo_module_diff_value_15, nx26514, nx26530, nx26542, 
         nx26544, nx26552, nx26566, camera_module_algo_module_prev_cont_value_15, 
         nx26580, camera_module_algo_module_prev_cont_value_14, nx26596, nx26604, 
         camera_module_algo_module_prev_cont_value_13, nx26612, 
         camera_module_algo_module_prev_cont_value_12, nx26628, nx26636, 
         camera_module_algo_module_prev_cont_value_11, nx26644, 
         camera_module_algo_module_prev_cont_value_10, nx26660, nx26668, 
         camera_module_algo_module_prev_cont_value_9, nx26676, 
         camera_module_algo_module_prev_cont_value_8, nx26692, nx26700, 
         camera_module_algo_module_prev_cont_value_7, nx26708, 
         camera_module_algo_module_prev_cont_value_6, nx26724, nx26732, 
         camera_module_algo_module_prev_cont_value_5, nx26740, 
         camera_module_algo_module_prev_cont_value_4, nx26756, nx26764, 
         camera_module_algo_module_prev_cont_value_3, nx26772, 
         camera_module_algo_module_prev_cont_value_2, nx26788, nx26796, 
         camera_module_algo_module_prev_cont_value_1, nx26804, 
         camera_module_algo_module_prev_cont_value_0, nx26820, nx26828, nx26844, 
         nx26860, nx26876, nx26892, nx26908, nx26924, nx26940, nx26956, 
         camera_module_algo_module_current_cont_value_16, 
         camera_module_algo_module_Addout_value_16, 
         camera_module_algo_module_diff_value_16, nx26970, nx26974, nx26984, 
         nx27002, nx27016, camera_module_algo_module_prev_cont_value_16, nx27030, 
         nx27038, camera_module_algo_module_failure_count_value_0, 
         camera_module_algo_module_modCU_current_state_14, nx27068, nx27084, 
         camera_module_algo_module_modCU_current_state_1, nx27106, nx27122, 
         nx27132, nx27156, nx27166, nx941, nx953, nx963, nx973, nx983, nx993, 
         nx1003, nx1013, nx1023, nx1033, nx1043, nx1053, nx1063, nx1073, nx1083, 
         nx1093, nx1103, nx1113, nx1123, nx1133, nx1143, nx1153, nx1163, nx1173, 
         nx1183, nx1193, nx1203, nx1213, nx1221, nx1233, nx1243, nx1253, nx1263, 
         nx1273, nx1283, nx1293, nx1303, nx1313, nx1323, nx1333, nx1343, nx1353, 
         nx1363, nx1373, nx1383, nx1393, nx1403, nx1413, nx1423, nx1433, nx1443, 
         nx1453, nx1463, nx1473, nx1483, nx1493, nx1503, nx1513, nx1523, nx1533, 
         nx1543, nx1553, nx1563, nx1573, nx1583, nx1593, nx1603, nx1613, nx1623, 
         nx1633, nx1643, nx1653, nx1663, nx1673, nx1683, nx1693, nx1703, nx1713, 
         nx1723, nx1733, nx1743, nx1753, nx1763, nx1773, nx1783, nx1793, nx1803, 
         nx1813, nx1823, nx1833, nx1843, nx1853, nx1863, nx1873, nx1883, nx1893, 
         nx1903, nx1913, nx1923, nx1933, nx1943, nx1953, nx1963, nx1973, nx1983, 
         nx1993, nx2003, nx2013, nx2023, nx2033, nx2043, nx2053, nx2063, nx2073, 
         nx2083, nx2093, nx2103, nx2113, nx2123, nx2133, nx2143, nx2153, nx2163, 
         nx2173, nx2183, nx2193, nx2203, nx2213, nx2223, nx2233, nx2243, nx2253, 
         nx2263, nx2273, nx2283, nx2293, nx2303, nx2313, nx2323, nx2333, nx2343, 
         nx2353, nx2363, nx2373, nx2383, nx2393, nx2403, nx2413, nx2423, nx2433, 
         nx2443, nx2453, nx2463, nx2473, nx2483, nx2493, nx2503, nx2513, nx2523, 
         nx2533, nx2543, nx2553, nx2563, nx2573, nx2583, nx2593, nx2603, nx2613, 
         nx2623, nx2633, nx2643, nx2653, nx2663, nx2673, nx2683, nx2693, nx2703, 
         nx2713, nx2723, nx2733, nx2743, nx2753, nx2763, nx2773, nx2783, nx2793, 
         nx2803, nx2813, nx2823, nx2833, nx2843, nx2853, nx2863, nx2873, nx2883, 
         nx2893, nx2903, nx2913, nx2923, nx2933, nx2943, nx2953, nx2963, nx2973, 
         nx2983, nx2993, nx3003, nx3013, nx3023, nx3033, nx3043, nx3053, nx3063, 
         nx3073, nx3083, nx3093, nx3103, nx3113, nx3123, nx3133, nx3143, nx3153, 
         nx3163, nx3173, nx3183, nx3193, nx3203, nx3213, nx3223, nx3233, nx3243, 
         nx3253, nx3263, nx3273, nx3283, nx3293, nx3303, nx3313, nx3323, nx3333, 
         nx3343, nx3353, nx3363, nx3373, nx3383, nx3393, nx3403, nx3413, nx3423, 
         nx3433, nx3443, nx3453, nx3463, nx3473, nx3483, nx3493, nx3503, nx3513, 
         nx3523, nx3533, nx3543, nx3553, nx3563, nx3573, nx3583, nx3593, nx3603, 
         nx3613, nx3623, nx3633, nx3643, nx3653, nx3663, nx3673, nx3683, nx3693, 
         nx3703, nx3713, nx3723, nx3733, nx3743, nx3753, nx3763, nx3773, nx3783, 
         nx3793, nx3803, nx3813, nx3823, nx3833, nx3843, nx3853, nx3863, nx3873, 
         nx3883, nx3893, nx3903, nx3913, nx3923, nx3933, nx3943, nx3953, nx3963, 
         nx3973, nx3983, nx3993, nx4003, nx4013, nx4023, nx4033, nx4043, nx4053, 
         nx4063, nx4073, nx4083, nx4093, nx4103, nx4113, nx4123, nx4133, nx4143, 
         nx4153, nx4163, nx4173, nx4183, nx4193, nx4203, nx4213, nx4223, nx4233, 
         nx4243, nx4253, nx4263, nx4273, nx4283, nx4293, nx4303, nx4313, nx4323, 
         nx4333, nx4343, nx4353, nx4363, nx4373, nx4383, nx4393, nx4403, nx4413, 
         nx4423, nx4433, nx4443, nx4453, nx4463, nx4473, nx4483, nx4493, nx4503, 
         nx4513, nx4523, nx4533, nx4543, nx4553, nx4563, nx4573, nx4583, nx4593, 
         nx4603, nx4613, nx4623, nx4633, nx4643, nx4653, nx4663, nx4673, nx4683, 
         nx4693, nx4703, nx4713, nx4723, nx4733, nx4743, nx4753, nx4763, nx4773, 
         nx4783, nx4793, nx4803, nx4813, nx4823, nx4833, nx4843, nx4853, nx4863, 
         nx4873, nx4883, nx4893, nx4903, nx4913, nx4923, nx4933, nx4943, nx4953, 
         nx4963, nx4973, nx4983, nx4993, nx5003, nx5013, nx5023, nx5033, nx5043, 
         nx5053, nx5063, nx5073, nx5083, nx5093, nx5103, nx5113, nx5123, nx5133, 
         nx5143, nx5153, nx5163, nx5173, nx5183, nx5193, nx5203, nx5213, nx5223, 
         nx5233, nx5243, nx5253, nx5263, nx5273, nx5283, nx5293, nx5303, nx5313, 
         nx5323, nx5333, nx5343, nx5353, nx5363, nx5373, nx5383, nx5393, nx5403, 
         nx5413, nx5423, nx5433, nx5443, nx5453, nx5463, nx5473, nx5483, nx5493, 
         nx5503, nx5513, nx5523, nx5533, nx5543, nx5553, nx5563, nx5573, nx5583, 
         nx5593, nx5603, nx5613, nx5623, nx5633, nx5643, nx5653, nx5663, nx5673, 
         nx5683, nx5693, nx5703, nx5713, nx5723, nx5733, nx5743, nx5753, nx5763, 
         nx5773, nx5783, nx5793, nx5803, nx5813, nx5823, nx5833, nx5843, nx5853, 
         nx5863, nx5873, nx5883, nx5893, nx5903, nx5913, nx5923, nx5933, nx5943, 
         nx5953, nx5963, nx5973, nx5983, nx5993, nx6003, nx6013, nx6023, nx6033, 
         nx6043, nx6053, nx6063, nx6073, nx6083, nx6093, nx6103, nx6113, nx6123, 
         nx6133, nx6143, nx6153, nx6163, nx6173, nx6183, nx6193, nx6203, nx6213, 
         nx6223, nx6233, nx6243, nx6253, nx6263, nx6273, nx6283, nx6293, nx6303, 
         nx6313, nx6323, nx6333, nx6343, nx6353, nx6363, nx6373, nx6383, nx6393, 
         nx6403, nx6413, nx6423, nx6433, nx6443, nx6453, nx6463, nx6473, nx6483, 
         nx6493, nx6503, nx6513, nx6523, nx6533, nx6543, nx6553, nx6563, nx6573, 
         nx6583, nx6593, nx6603, nx6613, nx6623, nx6633, nx6643, nx6653, nx6663, 
         nx6673, nx6683, nx6693, nx6703, nx6713, nx6723, nx6733, nx6743, nx6753, 
         nx6763, nx6773, nx6783, nx6793, nx6803, nx6813, nx6823, nx6833, nx6843, 
         nx6853, nx6863, nx6873, nx6883, nx6893, nx6903, nx6913, nx6923, nx6933, 
         nx6943, nx6953, nx6963, nx6973, nx6983, nx6993, nx7003, nx7013, nx7023, 
         nx7033, nx7043, nx7053, nx7063, nx7073, nx7083, nx7093, nx7103, nx7113, 
         nx7123, nx7133, nx7143, nx7153, nx7163, nx7173, nx7183, nx7193, nx7203, 
         nx7213, nx7223, nx7233, nx7243, nx7253, nx7263, nx7273, nx7283, nx7293, 
         nx7303, nx7313, nx7323, nx7333, nx7343, nx7353, nx7363, nx7373, nx7383, 
         nx7393, nx7403, nx7413, nx7423, nx7433, nx7443, nx7453, nx7463, nx7473, 
         nx7483, nx7493, nx7503, nx7513, nx7523, nx7533, nx7543, nx7553, nx7563, 
         nx7573, nx7583, nx7593, nx7603, nx7613, nx7623, nx7633, nx7643, nx7653, 
         nx7663, nx7673, nx7683, nx7693, nx7703, nx7713, nx7723, nx7733, nx7743, 
         nx7753, nx7763, nx7773, nx7783, nx7793, nx7803, nx7813, nx7823, nx7833, 
         nx7843, nx7853, nx7863, nx7873, nx7883, nx7893, nx7903, nx7913, nx7923, 
         nx7933, nx7943, nx7953, nx7963, nx7973, nx7983, nx7993, nx8003, nx8013, 
         nx8023, nx8033, nx8043, nx8053, nx8063, nx8073, nx8083, nx8093, nx8103, 
         nx8113, nx8123, nx8133, nx8143, nx8153, nx8163, nx8173, nx8183, nx8193, 
         nx8203, nx8213, nx8223, nx8233, nx8243, nx8253, nx8263, nx8273, nx8283, 
         nx8293, nx8303, nx8313, nx8323, nx8333, nx8343, nx8353, nx8363, nx8373, 
         nx8383, nx8393, nx8403, nx8413, nx8423, nx8433, nx8443, nx8453, nx8463, 
         nx8473, nx8483, nx8493, nx8503, nx8513, nx8523, nx8533, nx8543, nx8553, 
         nx8563, nx8573, nx8583, nx8593, nx8603, nx8613, nx8623, nx8633, nx8643, 
         nx8653, nx8663, nx8673, nx8683, nx8693, nx8703, nx8713, nx8723, nx8733, 
         nx8743, nx8753, nx8763, nx8773, nx8783, nx8793, nx8803, nx8813, nx8823, 
         nx8833, nx8843, nx8853, nx8863, nx8873, nx8883, nx8893, nx8903, nx8913, 
         nx8923, nx8933, nx8943, nx8953, nx8963, nx8973, nx8983, nx8993, nx9003, 
         nx9013, nx9023, nx9033, nx9043, nx9053, nx9063, nx9073, nx9083, nx9093, 
         nx9103, nx9113, nx9123, nx9133, nx9143, nx9153, nx9163, nx9173, nx9183, 
         nx9193, nx9203, nx9213, nx9223, nx9233, nx9243, nx9253, nx9263, nx9273, 
         nx9283, nx9293, nx9303, nx9313, nx9323, nx9333, nx9343, nx9353, nx9363, 
         nx9373, nx9383, nx9393, nx9403, nx9413, nx9423, nx9433, nx9443, nx9453, 
         nx9463, nx9473, nx9483, nx9493, nx9503, nx9513, nx9523, nx9533, nx9543, 
         nx9553, nx9563, nx9573, nx9583, nx9593, nx9603, nx9613, nx9623, nx9633, 
         nx9643, nx9653, nx9663, nx9673, nx9683, nx9693, nx9703, nx9713, nx9723, 
         nx9733, nx9743, nx9753, nx9763, nx9773, nx9783, nx9793, nx9803, nx9813, 
         nx9823, nx9833, nx9843, nx9853, nx9863, nx9873, nx9883, nx9893, nx9903, 
         nx9913, nx9923, nx9933, nx9943, nx9953, nx9963, nx9973, nx9983, nx9993, 
         nx10003, nx10013, nx10023, nx10033, nx10043, nx10053, nx10063, nx10073, 
         nx10083, nx10093, nx10103, nx10113, nx10123, nx10133, nx10143, nx10153, 
         nx10163, nx10173, nx10183, nx10193, nx10203, nx10213, nx10223, nx10233, 
         nx10243, nx10253, nx10263, nx10273, nx10283, nx10293, nx10303, nx10313, 
         nx10323, nx10333, nx10343, nx10353, nx10363, nx10373, nx10383, nx10393, 
         nx10403, nx10413, nx10423, nx10433, nx10443, nx10453, nx10463, nx10473, 
         nx10483, nx10493, nx10503, nx10513, nx10523, nx10533, nx10543, nx10553, 
         nx10563, nx10573, nx10583, nx10593, nx10603, nx10613, nx10623, nx10633, 
         nx10643, nx10653, nx10663, nx10673, nx10683, nx10693, nx10703, nx10713, 
         nx10723, nx10733, nx10743, nx10753, nx10763, nx10773, nx10783, nx10793, 
         nx10803, nx10813, nx10823, nx10833, nx10843, nx10853, nx10863, nx10873, 
         nx10883, nx10893, nx10903, nx10913, nx10923, nx10933, nx10943, nx10953, 
         nx10963, nx10973, nx10983, nx10993, nx11003, nx11013, nx11023, nx11033, 
         nx11043, nx11053, nx11063, nx11073, nx11083, nx11093, nx11103, nx11113, 
         nx11123, nx11133, nx11143, nx11153, nx11163, nx11173, nx11183, nx11193, 
         nx11203, nx11213, nx11223, nx11233, nx11243, nx11253, nx11263, nx11273, 
         nx11283, nx11293, nx11303, nx11313, nx11323, nx11333, nx11343, nx11353, 
         nx11363, nx11373, nx11383, nx11393, nx11403, nx11413, nx11423, nx11433, 
         nx11443, nx11453, nx11463, nx11473, nx11483, nx11493, nx11503, nx11513, 
         nx11523, nx11533, nx11543, nx11553, nx11563, nx11573, nx11583, nx11593, 
         nx11603, nx11613, nx11623, nx11633, nx11643, nx11653, nx11663, nx11673, 
         nx11683, nx11693, nx11703, nx11713, nx11723, nx11733, nx11743, nx11753, 
         nx11763, nx11773, nx11783, nx11793, nx11803, nx11813, nx11823, nx11833, 
         nx11843, nx11853, nx11863, nx11873, nx11883, nx11893, nx11903, nx11913, 
         nx11923, nx11933, nx11943, nx11953, nx11963, nx11973, nx11983, nx11993, 
         nx12003, nx12013, nx12023, nx12033, nx12043, nx12053, nx12063, nx12073, 
         nx12083, nx12093, nx12103, nx12113, nx12123, nx12133, nx12143, nx12153, 
         nx12163, nx12173, nx12183, nx12193, nx12203, nx12213, nx12223, nx12233, 
         nx12243, nx12253, nx12263, nx12273, nx12283, nx12293, nx12303, nx12313, 
         nx12323, nx12333, nx12343, nx12353, nx12363, nx12373, nx12383, nx12393, 
         nx12403, nx12413, nx12423, nx12433, nx12443, nx12453, nx12463, nx12473, 
         nx12483, nx12493, nx12503, nx12513, nx12523, nx12533, nx12543, nx12553, 
         nx12563, nx12573, nx12583, nx12593, nx12603, nx12613, nx12623, nx12633, 
         nx12643, nx12653, nx12663, nx12673, nx12683, nx12693, nx12703, nx12713, 
         nx12723, nx12733, nx12743, nx12753, nx12763, nx12773, nx12783, nx12793, 
         nx12803, nx12813, nx12823, nx12833, nx12843, nx12853, nx12863, nx12873, 
         nx12883, nx12893, nx12903, nx12913, nx12923, nx12933, nx12943, nx12953, 
         nx12963, nx12973, nx12983, nx12993, nx13003, nx13013, nx13023, nx13033, 
         nx13043, nx13053, nx13063, nx13073, nx13083, nx13093, nx13103, nx13113, 
         nx13123, nx13133, nx13143, nx13153, nx13163, nx13173, nx13183, nx13193, 
         nx13203, nx13213, nx13223, nx13233, nx13243, nx13253, nx13263, nx13273, 
         nx13283, nx13293, nx13303, nx13313, nx13323, nx13333, nx13343, nx13353, 
         nx13363, nx13373, nx13383, nx13393, nx13403, nx13413, nx13423, nx13433, 
         nx13443, nx13453, nx13463, nx13473, nx13483, nx13493, nx13503, nx13513, 
         nx13523, nx13533, nx13543, nx13553, nx13563, nx13573, nx13583, nx13593, 
         nx13603, nx13613, nx13623, nx13633, nx13643, nx13653, nx13663, nx13673, 
         nx13683, nx13693, nx13703, nx13713, nx13723, nx13733, nx13743, nx13753, 
         nx13763, nx13773, nx13783, nx13793, nx13803, nx13813, nx13823, nx13833, 
         nx13843, nx13853, nx13863, nx13873, nx13883, nx13893, nx13903, nx13913, 
         nx13923, nx13933, nx13943, nx13953, nx13963, nx13973, nx13983, nx13993, 
         nx14003, nx14013, nx14023, nx14033, nx14043, nx14053, nx14063, nx14073, 
         nx14083, nx14093, nx14103, nx14113, nx14123, nx14133, nx14143, nx14153, 
         nx14163, nx14173, nx14183, nx14193, nx14203, nx14213, nx14223, nx14233, 
         nx14243, nx14253, nx14263, nx14273, nx14283, nx14293, nx14303, nx14313, 
         nx14323, nx14333, nx14343, nx14353, nx14363, nx14373, nx14383, nx14393, 
         nx14403, nx14413, nx14423, nx14433, nx14443, nx14453, nx14463, nx14473, 
         nx14483, nx14493, nx14503, nx14513, nx14523, nx14533, nx14543, nx14553, 
         nx14563, nx14573, nx14583, nx14593, nx14603, nx14613, nx14623, nx14633, 
         nx14643, nx14653, nx14663, nx14673, nx14683, nx14693, nx14703, nx14713, 
         nx14723, nx14733, nx14743, nx14753, nx14763, nx14773, nx14783, nx14793, 
         nx14803, nx14813, nx14823, nx14833, nx14843, nx14853, nx14863, nx14873, 
         nx14883, nx14893, nx14903, nx14913, nx14923, nx14933, nx14943, nx14953, 
         nx14963, nx14973, nx14983, nx14993, nx15003, nx15013, nx15023, nx15033, 
         nx15043, nx15053, nx15063, nx15073, nx15083, nx15093, nx15103, nx15113, 
         nx15123, nx15133, nx15143, nx15153, nx15163, nx15173, nx15183, nx15193, 
         nx15203, nx15213, nx15223, nx15233, nx15243, nx15253, nx15263, nx15273, 
         nx15283, nx15293, nx15303, nx15313, nx15323, nx15333, nx15343, nx15353, 
         nx15363, nx15373, nx15383, nx15393, nx15403, nx15413, nx15423, nx15433, 
         nx15443, nx15453, nx15463, nx15473, nx15483, nx15493, nx15503, nx15513, 
         nx15523, nx15533, nx15543, nx15553, nx15563, nx15573, nx15583, nx15593, 
         nx15603, nx15613, nx15623, nx15633, nx15643, nx15653, nx15663, nx15673, 
         nx15683, nx15693, nx15703, nx15713, nx15723, nx15733, nx15743, nx15753, 
         nx15763, nx15773, nx15783, nx15793, nx15803, nx15813, nx15823, nx15833, 
         nx15843, nx15853, nx15863, nx15873, nx15883, nx15893, nx15903, nx15913, 
         nx15923, nx15933, nx15943, nx15953, nx15963, nx15973, nx15983, nx15993, 
         nx16003, nx16013, nx16023, nx16033, nx16043, nx16053, nx16063, nx16073, 
         nx16083, nx16093, nx16103, nx16113, nx16123, nx16133, nx16143, nx16153, 
         nx16163, nx16173, nx16183, nx16193, nx16203, nx16213, nx16223, nx16233, 
         nx16243, nx16253, nx16263, nx16273, nx16283, nx16293, nx16303, nx16313, 
         nx16323, nx16333, nx16343, nx16353, nx16363, nx16373, nx16383, nx16393, 
         nx16403, nx16413, nx16423, nx16433, nx16443, nx16453, nx16463, nx16473, 
         nx16483, nx16493, nx16503, nx16513, nx16523, nx16533, nx16543, nx16553, 
         nx16563, nx16573, nx16583, nx16593, nx16603, nx16613, nx16623, nx16633, 
         nx16643, nx16653, nx16663, nx16673, nx16683, nx16693, nx16703, nx16713, 
         nx16723, nx16733, nx16743, nx16753, nx16763, nx16773, nx16783, nx16793, 
         nx16803, nx16813, nx16823, nx16833, nx16843, nx16853, nx16863, nx16873, 
         nx16883, nx16893, nx16903, nx16913, nx16923, nx16933, nx16943, nx16953, 
         nx16963, nx16973, nx16983, nx16993, nx17003, nx17013, nx17023, nx17033, 
         nx17043, nx17053, nx17063, nx17073, nx17083, nx17093, nx17103, nx17113, 
         nx17123, nx17133, nx17143, nx17153, nx17163, nx17173, nx17183, nx17193, 
         nx17203, nx17213, nx17223, nx17233, nx17243, nx17253, nx17263, nx17273, 
         nx17283, nx17293, nx17303, nx17313, nx17323, nx17333, nx17343, nx17353, 
         nx17363, nx17373, nx17383, nx17393, nx17403, nx17413, nx17423, nx17433, 
         nx17443, nx17453, nx17463, nx17473, nx17483, nx17493, nx17503, nx17513, 
         nx17523, nx17533, nx17543, nx17553, nx17563, nx17573, nx17583, nx17593, 
         nx17603, nx17613, nx17623, nx17633, nx17643, nx17653, nx17663, nx17673, 
         nx17683, nx17693, nx17703, nx17713, nx17723, nx17733, nx17743, nx17753, 
         nx17763, nx17773, nx17783, nx17793, nx17803, nx17813, nx17823, nx17833, 
         nx17843, nx17853, nx17863, nx17873, nx17883, nx17893, nx17903, nx17913, 
         nx17923, nx17933, nx17943, nx17953, nx17963, nx17973, nx17983, nx17993, 
         nx18003, nx18013, nx18023, nx18033, nx18043, nx18053, nx18063, nx18073, 
         nx18083, nx18093, nx18103, nx18113, nx18123, nx18133, nx18143, nx18153, 
         nx18163, nx18173, nx18183, nx18193, nx18203, nx18213, nx18223, nx18233, 
         nx18243, nx18253, nx18263, nx18273, nx18283, nx18293, nx18303, nx18313, 
         nx18323, nx18333, nx18343, nx18353, nx18363, nx18373, nx18383, nx18393, 
         nx18403, nx18413, nx18423, nx18433, nx18443, nx18453, nx18463, nx18473, 
         nx18483, nx18493, nx18503, nx18513, nx18523, nx18533, nx18543, nx18553, 
         nx18563, nx18573, nx18583, nx18593, nx18603, nx18613, nx18623, nx18633, 
         nx18643, nx18653, nx18663, nx18673, nx18683, nx18693, nx18703, nx18713, 
         nx18723, nx18733, nx18743, nx18753, nx18763, nx18773, nx18783, nx18793, 
         nx18803, nx18813, nx18823, nx18833, nx18843, nx18853, nx18863, nx18873, 
         nx18883, nx18893, nx18903, nx18913, nx18923, nx18933, nx18943, nx18953, 
         nx18963, nx18973, nx18983, nx18993, nx19003, nx19013, nx19023, nx19033, 
         nx19043, nx19053, nx19063, nx19073, nx19083, nx19093, nx19103, nx19113, 
         nx19123, nx19133, nx19143, nx19153, nx19163, nx19173, nx19183, nx19193, 
         nx19203, nx19213, nx19223, nx19233, nx19243, nx19253, nx19263, nx19273, 
         nx19283, nx19293, nx19303, nx19313, nx19323, nx19333, nx19343, nx19353, 
         nx19363, nx19373, nx19383, nx19393, nx19403, nx19413, nx19423, nx19433, 
         nx19443, nx19453, nx19463, nx19473, nx19483, nx19493, nx19503, nx19513, 
         nx19523, nx19533, nx19543, nx19553, nx19563, nx19573, nx19583, nx19593, 
         nx19603, nx19613, nx19623, nx19633, nx19643, nx19653, nx19663, nx19673, 
         nx19683, nx19693, nx19703, nx19713, nx19723, nx19733, nx19743, nx19753, 
         nx19763, nx19773, nx19783, nx19793, nx19803, nx19813, nx19823, nx19833, 
         nx19843, nx19853, nx19863, nx19873, nx19883, nx19893, nx19903, nx19913, 
         nx19923, nx19933, nx19943, nx19953, nx19963, nx19973, nx19983, nx19993, 
         nx20003, nx20013, nx20023, nx20033, nx20043, nx20053, nx20063, nx20073, 
         nx20083, nx20093, nx20103, nx20113, nx20123, nx20133, nx20143, nx20153, 
         nx20163, nx20173, nx20183, nx20193, nx20203, nx20213, nx20223, nx20233, 
         nx20243, nx20253, nx20263, nx20273, nx20283, nx20293, nx20303, nx20313, 
         nx20323, nx20333, nx20343, nx20353, nx20363, nx20373, nx20383, nx20393, 
         nx20403, nx20413, nx20423, nx20433, nx20443, nx20453, nx20463, nx20473, 
         nx20483, nx20493, nx20503, nx20513, nx20523, nx20533, nx20543, nx20553, 
         nx20563, nx20573, nx20583, nx20593, nx20603, nx20613, nx20623, nx20633, 
         nx20643, nx20653, nx20663, nx20673, nx20683, nx20693, nx20703, nx20713, 
         nx20723, nx20733, nx20743, nx20753, nx20763, nx20773, nx20783, nx20793, 
         nx20803, nx20813, nx20823, nx20833, nx20843, nx20853, nx20863, nx20873, 
         nx20883, nx20893, nx20903, nx20913, nx20923, nx20933, nx20943, nx20953, 
         nx20963, nx20973, nx20983, nx20993, nx21003, nx21013, nx21023, nx21033, 
         nx21043, nx21053, nx21063, nx21073, nx21083, nx21093, nx21103, nx21113, 
         nx21123, nx21133, nx21143, nx21153, nx21163, nx21173, nx21183, nx21193, 
         nx21203, nx21213, nx21223, nx21233, nx21243, nx21253, nx21263, nx21273, 
         nx21283, nx21293, nx21303, nx21313, nx21323, nx21333, nx21343, nx21353, 
         nx21363, nx21373, nx21383, nx21393, nx21403, nx21413, nx21423, nx21433, 
         nx21443, nx21453, nx21463, nx21473, nx21483, nx21493, nx21503, nx21513, 
         nx21523, nx21533, nx21543, nx21553, nx21563, nx21573, nx21583, nx21593, 
         nx21603, nx21613, nx21623, nx21633, nx21643, nx21653, nx21663, nx21673, 
         nx21683, nx21693, nx21703, nx21713, nx21723, nx21733, nx21743, nx21753, 
         nx21763, nx21773, nx21783, nx21793, nx21803, nx21813, nx21823, nx21833, 
         nx21843, nx21853, nx21863, nx21873, nx21883, nx21893, nx21903, nx21913, 
         nx21923, nx21933, nx21943, nx21953, nx21963, nx21973, nx21983, nx21993, 
         nx22003, nx22013, nx22023, nx22033, nx22043, nx22053, nx22063, nx22073, 
         nx22083, nx22093, nx22103, nx22113, nx22123, nx22133, nx22143, nx22153, 
         nx22163, nx22173, nx22183, nx22193, nx22203, nx22213, nx22223, nx22233, 
         nx22243, nx22253, nx22263, nx22273, nx22283, nx22293, nx22303, nx22313, 
         nx22323, nx22333, nx22343, nx22353, nx22363, nx22373, nx22383, nx22393, 
         nx22403, nx22413, nx22423, nx22433, nx22443, nx22453, nx22463, nx22473, 
         nx22481, nx22493, nx22503, nx22513, nx22523, nx22533, nx22543, nx22549, 
         nx22565, nx22568, nx22575, nx22577, nx22579, nx22585, nx22587, nx22595, 
         nx22597, nx22601, nx22605, nx22611, nx22613, nx22627, nx22631, nx22645, 
         nx22651, nx22653, nx22665, nx22669, nx22677, nx22679, nx22681, nx22685, 
         nx22689, nx22693, nx22699, nx22701, nx22705, nx22709, nx22719, nx22727, 
         nx22739, nx22749, nx22753, nx22757, nx22761, nx22766, nx22771, nx22773, 
         nx22775, nx22777, nx22779, nx22787, nx22791, nx22795, nx22801, nx22805, 
         nx22811, nx22815, nx22821, nx22823, nx22825, nx22827, nx22831, nx22835, 
         nx22837, nx22839, nx22841, nx22844, nx22846, nx22849, nx22851, nx22871, 
         nx22874, nx22887, nx22891, nx22897, nx22907, nx22912, nx22915, nx22923, 
         nx22931, nx22935, nx22943, nx22945, nx22951, nx22953, nx22961, nx22963, 
         nx22968, nx22973, nx22979, nx22981, nx22987, nx22989, nx22993, nx22997, 
         nx23003, nx23005, nx23006, nx23011, nx23012, nx23016, nx23019, nx23021, 
         nx23026, nx23033, nx23051, nx23053, nx23055, nx23059, nx23067, nx23069, 
         nx23071, nx23073, nx23079, nx23084, nx23087, nx23091, nx23100, nx23102, 
         nx23105, nx23111, nx23113, nx23117, nx23119, nx23130, nx23138, nx23145, 
         nx23157, nx23165, nx23172, nx23189, nx23211, nx23218, nx23236, nx23256, 
         nx23267, nx23279, nx23282, nx23290, nx23298, nx23302, nx23305, nx23314, 
         nx23324, nx23337, nx23349, nx23361, nx23372, nx23385, nx23400, nx23413, 
         nx23417, nx23423, nx23433, nx23446, nx23458, nx23469, nx23482, nx23495, 
         nx23506, nx23520, nx23523, nx23529, nx23537, nx23549, nx23562, nx23574, 
         nx23587, nx23599, nx23610, nx23627, nx23630, nx23639, nx23648, nx23660, 
         nx23670, nx23683, nx23695, nx23706, nx23719, nx23733, nx23736, nx23748, 
         nx23761, nx23772, nx23785, nx23797, nx23811, nx23822, nx23835, nx23839, 
         nx23852, nx23863, nx23875, nx23889, nx23900, nx23913, nx23925, nx23938, 
         nx23941, nx23954, nx23966, nx23977, nx23989, nx24001, nx24012, nx24024, 
         nx24041, nx24045, nx24053, nx24060, nx24073, nx24084, nx24097, nx24109, 
         nx24120, nx24133, nx24146, nx24149, nx24162, nx24174, nx24184, nx24197, 
         nx24209, nx24222, nx24235, nx24248, nx24251, nx24264, nx24276, nx24286, 
         nx24300, nx24313, nx24324, nx24336, nx24349, nx24353, nx24364, nx24379, 
         nx24390, nx24403, nx24415, nx24428, nx24440, nx24455, nx24459, nx24463, 
         nx24473, nx24477, nx24481, nx24487, nx24490, nx24495, nx24500, nx24503, 
         nx24508, nx24513, nx24517, nx24521, nx24526, nx24529, nx24535, nx24541, 
         nx24544, nx24548, nx24554, nx24557, nx24563, nx24569, nx24572, nx24575, 
         nx24581, nx24589, nx24592, nx24597, nx24602, nx24605, nx24610, nx24615, 
         nx24619, nx24624, nx24629, nx24633, nx24637, nx24642, nx24645, nx24650, 
         nx24655, nx24659, nx24663, nx24669, nx24672, nx24677, nx24682, nx24686, 
         nx24689, nx24693, nx24703, nx24707, nx24712, nx24717, nx24720, nx24725, 
         nx24730, nx24733, nx24738, nx24743, nx24747, nx24751, nx24757, nx24760, 
         nx24765, nx24770, nx24774, nx24778, nx24785, nx24788, nx24792, nx24798, 
         nx24801, nx24805, nx24809, nx24811, nx24816, nx24819, nx24825, nx24830, 
         nx24834, nx24838, nx24845, nx24848, nx24853, nx24859, nx24863, nx24869, 
         nx24874, nx24877, nx24882, nx24887, nx24890, nx24894, nx24900, nx24903, 
         nx24909, nx24914, nx24918, nx24921, nx24925, nx24930, nx24933, nx24935, 
         nx24939, nx24945, nx24947, nx24951, nx24954, nx24960, nx24979, nx24983, 
         nx24997, nx25001, nx25009, nx25017, nx25027, nx25039, nx25047, nx25056, 
         nx25065, nx25074, nx25077, nx25085, nx25094, nx25103, nx25113, nx25122, 
         nx25131, nx25140, nx25149, nx25153, nx25162, nx25172, nx25181, nx25191, 
         nx25201, nx25209, nx25218, nx25227, nx25231, nx25241, nx25251, nx25261, 
         nx25271, nx25281, nx25291, nx25301, nx25311, nx25315, nx25324, nx25334, 
         nx25343, nx25353, nx25365, nx25376, nx25386, nx25397, nx25401, nx25413, 
         nx25425, nx25437, nx25449, nx25459, nx25469, nx25480, nx25489, nx25493, 
         nx25502, nx25515, nx25525, nx25536, nx25549, nx25559, nx25568, nx25576, 
         nx25581, nx25593, nx25604, nx25613, nx25625, nx25634, nx25644, nx25655, 
         nx25667, nx25671, nx25681, nx25691, nx25702, nx25711, nx25721, nx25733, 
         nx25744, nx25754, nx25757, nx25768, nx25778, nx25787, nx25797, nx25809, 
         nx25821, nx25831, nx25842, nx25845, nx25855, nx25864, nx25872, nx25885, 
         nx25895, nx25905, nx25916, nx25926, nx25929, nx25938, nx25946, nx25959, 
         nx25969, nx25979, nx25990, nx26000, nx26009, nx26013, nx26023, nx26034, 
         nx26045, nx26055, nx26067, nx26077, nx26086, nx26094, nx26099, nx26111, 
         nx26122, nx26131, nx26143, nx26152, nx26162, nx26173, nx26185, nx26189, 
         nx26199, nx26209, nx26220, nx26229, nx26239, nx26251, nx26262, nx26272, 
         nx26275, nx26286, nx26296, nx26305, nx26315, nx26327, nx26339, nx26349, 
         nx26363, nx26370, nx26372, nx26375, nx26379, nx26385, nx26411, nx26415, 
         nx26429, nx26435, nx26444, nx26453, nx26463, nx26475, nx26487, nx26497, 
         nx26508, nx26521, nx26525, nx26536, nx26545, nx26554, nx26563, nx26573, 
         nx26582, nx26590, nx26600, nx26603, nx26614, nx26622, nx26632, nx26643, 
         nx26653, nx26662, nx26670, nx26680, nx26683, nx26694, nx26702, nx26712, 
         nx26723, nx26733, nx26742, nx26750, nx26761, nx26765, nx26774, nx26782, 
         nx26792, nx26803, nx26813, nx26822, nx26831, nx26843, nx26847, nx26859, 
         nx26871, nx26883, nx26895, nx26907, nx26919, nx26931, nx26943, nx26947, 
         nx26959, nx26971, nx26983, nx26993, nx27004, nx27013, nx27023, nx27032, 
         nx27035, nx27045, nx27054, nx27065, nx27076, nx27088, nx27097, nx27105, 
         nx27115, nx27119, nx27131, nx27142, nx27152, nx27163, nx27173, nx27181, 
         nx27189, nx27197, nx27200, nx27208, nx27216, nx27224, nx27233, nx27241, 
         nx27249, nx27257, nx27265, nx27268, nx27276, nx27284, nx27292, nx27301, 
         nx27309, nx27317, nx27325, nx27333, nx27336, nx27344, nx27352, nx27360, 
         nx27369, nx27377, nx27385, nx27393, nx27402, nx27405, nx27413, nx27421, 
         nx27429, nx27438, nx27446, nx27454, nx27462, nx27470, nx27473, nx27481, 
         nx27489, nx27497, nx27506, nx27514, nx27522, nx27530, nx27538, nx27541, 
         nx27549, nx27557, nx27565, nx27574, nx27582, nx27590, nx27598, nx27606, 
         nx27609, nx27617, nx27625, nx27633, nx27642, nx27650, nx27658, nx27666, 
         nx27676, nx27681, nx27683, nx27686, nx27689, nx27694, nx27710, nx27713, 
         nx27724, nx27728, nx27735, nx27743, nx27751, nx27760, nx27768, nx27776, 
         nx27784, nx27792, nx27795, nx27803, nx27811, nx27819, nx27828, nx27836, 
         nx27844, nx27852, nx27860, nx27863, nx27871, nx27879, nx27887, nx27896, 
         nx27904, nx27912, nx27920, nx27928, nx27931, nx27939, nx27947, nx27955, 
         nx27964, nx27972, nx27980, nx27988, nx27997, nx28000, nx28008, nx28016, 
         nx28024, nx28033, nx28041, nx28049, nx28057, nx28065, nx28068, nx28076, 
         nx28084, nx28092, nx28101, nx28109, nx28117, nx28125, nx28133, nx28136, 
         nx28144, nx28152, nx28160, nx28169, nx28177, nx28185, nx28193, nx28201, 
         nx28204, nx28212, nx28220, nx28228, nx28237, nx28245, nx28253, nx28261, 
         nx28270, nx28273, nx28281, nx28289, nx28297, nx28306, nx28314, nx28322, 
         nx28330, nx28338, nx28341, nx28349, nx28357, nx28365, nx28374, nx28382, 
         nx28390, nx28398, nx28406, nx28409, nx28417, nx28425, nx28433, nx28442, 
         nx28450, nx28458, nx28466, nx28474, nx28477, nx28485, nx28493, nx28501, 
         nx28510, nx28518, nx28526, nx28534, nx28543, nx28546, nx28554, nx28562, 
         nx28570, nx28579, nx28587, nx28595, nx28603, nx28611, nx28614, nx28622, 
         nx28630, nx28638, nx28647, nx28655, nx28663, nx28671, nx28679, nx28682, 
         nx28690, nx28698, nx28706, nx28715, nx28723, nx28731, nx28739, nx28747, 
         nx28750, nx28758, nx28766, nx28774, nx28783, nx28791, nx28799, nx28807, 
         nx28817, nx28822, nx28824, nx28827, nx28830, nx28835, nx28851, nx28854, 
         nx28865, nx28869, nx28876, nx28884, nx28892, nx28901, nx28909, nx28917, 
         nx28925, nx28933, nx28936, nx28944, nx28952, nx28960, nx28969, nx28977, 
         nx28985, nx28993, nx29001, nx29004, nx29012, nx29020, nx29028, nx29037, 
         nx29045, nx29053, nx29061, nx29069, nx29072, nx29080, nx29088, nx29096, 
         nx29105, nx29113, nx29121, nx29129, nx29138, nx29141, nx29149, nx29157, 
         nx29165, nx29174, nx29182, nx29190, nx29198, nx29206, nx29209, nx29217, 
         nx29225, nx29233, nx29242, nx29250, nx29258, nx29266, nx29274, nx29277, 
         nx29285, nx29293, nx29301, nx29310, nx29318, nx29326, nx29334, nx29342, 
         nx29345, nx29353, nx29361, nx29369, nx29378, nx29386, nx29394, nx29402, 
         nx29411, nx29414, nx29422, nx29430, nx29438, nx29447, nx29455, nx29463, 
         nx29471, nx29479, nx29482, nx29490, nx29498, nx29506, nx29515, nx29523, 
         nx29531, nx29539, nx29547, nx29550, nx29558, nx29566, nx29574, nx29583, 
         nx29591, nx29599, nx29607, nx29615, nx29618, nx29626, nx29634, nx29642, 
         nx29651, nx29659, nx29667, nx29675, nx29684, nx29687, nx29695, nx29703, 
         nx29711, nx29720, nx29728, nx29736, nx29744, nx29752, nx29755, nx29763, 
         nx29771, nx29779, nx29788, nx29796, nx29804, nx29812, nx29820, nx29823, 
         nx29831, nx29839, nx29847, nx29856, nx29864, nx29872, nx29880, nx29888, 
         nx29891, nx29899, nx29907, nx29915, nx29924, nx29932, nx29940, nx29948, 
         nx29956, nx29959, nx29964, nx29966, nx29969, nx29972, nx29977, nx29993, 
         nx29996, nx30007, nx30011, nx30018, nx30026, nx30034, nx30043, nx30051, 
         nx30059, nx30067, nx30075, nx30078, nx30086, nx30094, nx30102, nx30111, 
         nx30119, nx30127, nx30135, nx30143, nx30146, nx30154, nx30162, nx30170, 
         nx30179, nx30187, nx30195, nx30203, nx30211, nx30214, nx30222, nx30230, 
         nx30238, nx30247, nx30255, nx30263, nx30271, nx30280, nx30283, nx30291, 
         nx30299, nx30307, nx30316, nx30324, nx30332, nx30340, nx30348, nx30351, 
         nx30359, nx30367, nx30375, nx30384, nx30392, nx30400, nx30408, nx30416, 
         nx30419, nx30427, nx30435, nx30443, nx30452, nx30460, nx30468, nx30476, 
         nx30484, nx30487, nx30495, nx30503, nx30511, nx30520, nx30528, nx30536, 
         nx30544, nx30553, nx30556, nx30564, nx30572, nx30580, nx30589, nx30597, 
         nx30605, nx30613, nx30621, nx30624, nx30632, nx30640, nx30648, nx30657, 
         nx30665, nx30673, nx30681, nx30689, nx30692, nx30700, nx30708, nx30716, 
         nx30725, nx30733, nx30741, nx30749, nx30757, nx30760, nx30768, nx30776, 
         nx30784, nx30793, nx30801, nx30809, nx30817, nx30826, nx30829, nx30837, 
         nx30845, nx30853, nx30862, nx30870, nx30878, nx30886, nx30894, nx30897, 
         nx30905, nx30913, nx30921, nx30930, nx30938, nx30946, nx30954, nx30962, 
         nx30965, nx30973, nx30981, nx30989, nx30998, nx31006, nx31014, nx31022, 
         nx31030, nx31033, nx31041, nx31049, nx31057, nx31066, nx31074, nx31082, 
         nx31090, nx31098, nx31101, nx31106, nx31108, nx31111, nx31114, nx31119, 
         nx31135, nx31138, nx31149, nx31153, nx31160, nx31168, nx31176, nx31185, 
         nx31193, nx31201, nx31209, nx31217, nx31220, nx31228, nx31236, nx31244, 
         nx31253, nx31261, nx31269, nx31277, nx31285, nx31288, nx31296, nx31304, 
         nx31312, nx31321, nx31329, nx31337, nx31345, nx31353, nx31356, nx31364, 
         nx31372, nx31380, nx31389, nx31397, nx31405, nx31413, nx31422, nx31425, 
         nx31433, nx31441, nx31449, nx31458, nx31466, nx31474, nx31482, nx31490, 
         nx31493, nx31501, nx31509, nx31517, nx31526, nx31534, nx31542, nx31550, 
         nx31558, nx31561, nx31569, nx31577, nx31585, nx31594, nx31602, nx31610, 
         nx31618, nx31626, nx31629, nx31637, nx31645, nx31653, nx31662, nx31670, 
         nx31678, nx31686, nx31695, nx31698, nx31706, nx31714, nx31722, nx31731, 
         nx31739, nx31747, nx31755, nx31763, nx31766, nx31774, nx31782, nx31790, 
         nx31799, nx31807, nx31815, nx31823, nx31831, nx31834, nx31842, nx31850, 
         nx31858, nx31867, nx31875, nx31883, nx31891, nx31899, nx31902, nx31910, 
         nx31918, nx31926, nx31935, nx31943, nx31951, nx31959, nx31968, nx31971, 
         nx31979, nx31987, nx31995, nx32004, nx32012, nx32020, nx32028, nx32036, 
         nx32039, nx32047, nx32055, nx32063, nx32072, nx32080, nx32088, nx32096, 
         nx32104, nx32107, nx32115, nx32123, nx32131, nx32140, nx32148, nx32156, 
         nx32164, nx32172, nx32175, nx32183, nx32191, nx32199, nx32208, nx32216, 
         nx32224, nx32232, nx32240, nx32243, nx32248, nx32250, nx32253, nx32256, 
         nx32261, nx32277, nx32280, nx32291, nx32295, nx32302, nx32310, nx32318, 
         nx32327, nx32335, nx32343, nx32351, nx32359, nx32362, nx32370, nx32378, 
         nx32386, nx32395, nx32403, nx32411, nx32419, nx32427, nx32430, nx32438, 
         nx32446, nx32454, nx32463, nx32471, nx32479, nx32487, nx32495, nx32498, 
         nx32506, nx32514, nx32522, nx32531, nx32539, nx32547, nx32555, nx32564, 
         nx32567, nx32575, nx32583, nx32591, nx32600, nx32608, nx32616, nx32624, 
         nx32632, nx32635, nx32643, nx32651, nx32659, nx32668, nx32676, nx32684, 
         nx32692, nx32700, nx32703, nx32711, nx32719, nx32727, nx32736, nx32744, 
         nx32752, nx32760, nx32768, nx32771, nx32779, nx32787, nx32795, nx32804, 
         nx32812, nx32820, nx32828, nx32837, nx32840, nx32848, nx32856, nx32864, 
         nx32873, nx32881, nx32889, nx32897, nx32905, nx32908, nx32916, nx32924, 
         nx32932, nx32941, nx32949, nx32957, nx32965, nx32973, nx32976, nx32984, 
         nx32992, nx33000, nx33009, nx33017, nx33025, nx33033, nx33041, nx33044, 
         nx33052, nx33060, nx33068, nx33077, nx33085, nx33093, nx33101, nx33110, 
         nx33113, nx33121, nx33129, nx33137, nx33146, nx33154, nx33162, nx33170, 
         nx33178, nx33181, nx33189, nx33197, nx33205, nx33214, nx33222, nx33230, 
         nx33238, nx33246, nx33249, nx33257, nx33265, nx33273, nx33282, nx33290, 
         nx33298, nx33306, nx33314, nx33317, nx33325, nx33333, nx33341, nx33350, 
         nx33358, nx33366, nx33374, nx33382, nx33384, nx33386, nx33388, nx33391, 
         nx33393, nx33396, nx33398, nx33401, nx33403, nx33405, nx33408, nx33410, 
         nx33412, nx33415, nx33419, nx33423, nx33425, nx33427, nx33429, nx33433, 
         nx33435, nx33437, nx33439, nx33444, nx33446, nx33451, nx33453, nx33458, 
         nx33460, nx33465, nx33467, nx33472, nx33474, nx33485, nx33489, nx33491, 
         nx33494, nx33504, nx33508, nx33510, nx33513, nx33523, nx33529, nx33540, 
         nx33546, nx33557, nx33563, nx33574, nx33580, nx33591, nx33608, nx33609, 
         nx33615, nx33616, nx33619, nx33621, nx33629, nx33632, nx33638, nx33639, 
         nx33642, nx33644, nx33652, nx33655, nx33661, nx33662, nx33665, nx33667, 
         nx33675, nx33678, nx33684, nx33685, nx33688, nx33690, nx33698, nx33701, 
         nx33707, nx33708, nx33711, nx33713, nx33721, nx33724, nx33727, nx33729, 
         nx33732, nx33734, nx33737, nx33739, nx33747, nx33750, nx33753, nx33755, 
         nx33758, nx33760, nx33763, nx33765, nx33773, nx33776, nx33779, nx33781, 
         nx33784, nx33790, nx33794, nx33796, nx33799, nx33801, nx33803, nx33805, 
         nx33807, nx33810, nx33816, nx33818, nx33825, nx33832, nx33834, nx33841, 
         nx33848, nx33850, nx33857, nx33864, nx33866, nx33873, nx33880, nx33882, 
         nx33889, nx33896, nx33898, nx33905, nx33912, nx33914, nx33921, nx33928, 
         nx33930, nx33943, nx33945, nx33948, nx33953, nx33958, nx33961, nx34003, 
         nx34005, nx34007, nx34010, nx34018, nx34027, nx34036, nx34038, nx34040, 
         nx34042, nx34066, nx34068, nx34070, nx34072, nx34074, nx34076, nx34080, 
         nx34082, nx34084, nx34086, nx34090, nx34092, nx34094, nx34096, nx34098, 
         nx34100, nx34102, nx34104, nx34106, nx34108, nx34110, nx34112, nx34118, 
         nx34120, nx34122, nx34124, nx34130, nx34132, nx34138, nx34140, nx34142, 
         nx34150, nx34164, nx34166, nx34168, nx34170, nx34172, nx34174, nx34176, 
         nx34178, nx34180, nx34182, nx34184, nx34186, nx34188, nx34190, nx34192, 
         nx34194, nx34196, nx34198, nx34200, nx34202, nx34204, nx34206, nx34208, 
         nx34210, nx34212, nx34214, nx34216, nx34218, nx34220, nx34222, nx34224, 
         nx34226, nx34228, nx34230, nx34232, nx34234, nx34236, nx34304, nx34306, 
         nx34308, nx34310, nx34312, nx34314, nx34316, nx34318, nx34320, nx34322, 
         nx34324, nx34326, nx34328, nx34330, nx34332, nx34334, nx34336, nx34338, 
         nx34340, nx34342, nx34344, nx34346, nx34348, nx34350, nx34352, nx34354, 
         nx34356, nx34358, nx34360, nx34362, nx34364, nx34366, nx34374, nx34376, 
         nx34378, nx34380, nx34382, nx34384, nx34386, nx34388, nx34390, nx34392, 
         nx34394, nx34396, nx34398, nx34400, nx34402, nx34404, nx34406, nx34408, 
         nx34410, nx34412, nx34414, nx34416, nx34418, nx34420, nx34422, nx34424, 
         nx34426, nx34428, nx34430, nx34432, nx34434, nx34436, nx34444, nx34446, 
         nx34448, nx34450, nx34452, nx34454, nx34456, nx34458, nx34460, nx34462, 
         nx34464, nx34466, nx34468, nx34470, nx34472, nx34474, nx34476, nx34478, 
         nx34480, nx34482, nx34484, nx34486, nx34488, nx34490, nx34492, nx34494, 
         nx34496, nx34498, nx34500, nx34502, nx34504, nx34506, nx34514, nx34516, 
         nx34518, nx34520, nx34522, nx34524, nx34526, nx34528, nx34530, nx34532, 
         nx34534, nx34536, nx34538, nx34540, nx34542, nx34544, nx34546, nx34548, 
         nx34550, nx34552, nx34554, nx34556, nx34558, nx34560, nx34562, nx34564, 
         nx34566, nx34568, nx34570, nx34572, nx34574, nx34576, nx34584, nx34586, 
         nx34588, nx34590, nx34592, nx34594, nx34596, nx34598, nx34600, nx34602, 
         nx34604, nx34606, nx34608, nx34610, nx34612, nx34614, nx34616, nx34618, 
         nx34620, nx34622, nx34624, nx34626, nx34628, nx34630, nx34632, nx34634, 
         nx34636, nx34638, nx34640, nx34642, nx34644, nx34646, nx34654, nx34656, 
         nx34658, nx34660, nx34662, nx34664, nx34666, nx34668, nx34670, nx34672, 
         nx34674, nx34676, nx34678, nx34680, nx34682, nx34684, nx34686, nx34688, 
         nx34690, nx34692, nx34694, nx34696, nx34698, nx34700, nx34702, nx34704, 
         nx34706, nx34708, nx34710, nx34712, nx34714, nx34716, nx34724, nx34726, 
         nx34728, nx34730, nx34732, nx34734, nx34736, nx34738, nx34740, nx34742, 
         nx34744, nx34746, nx34748, nx34750, nx34752, nx34754, nx34756, nx34758, 
         nx34760, nx34762, nx34764, nx34766, nx34768, nx34770, nx34772, nx34774, 
         nx34776, nx34778, nx34780, nx34782, nx34784, nx34786, nx34794, nx34796, 
         nx34798, nx34800, nx34802, nx34804, nx34806, nx34808, nx34810, nx34812, 
         nx34814, nx34816, nx34818, nx34820, nx34822, nx34824, nx34826, nx34828, 
         nx34830, nx34832, nx34834, nx34836, nx34838, nx34840, nx34842, nx34844, 
         nx34846, nx34848, nx34850, nx34852, nx34854, nx34856, nx34864, nx34866, 
         nx34868, nx34870, nx34872, nx34874, nx34876, nx34878, nx34880, nx34882, 
         nx34884, nx34886, nx34888, nx34890, nx34892, nx34894, nx34896, nx34898, 
         nx34900, nx34902, nx34904, nx34906, nx34908, nx34910, nx34912, nx34914, 
         nx34916, nx34918, nx34920, nx34922, nx34924, nx34926, nx34934, nx34936, 
         nx34938, nx34940, nx34942, nx34944, nx34946, nx34948, nx34950, nx34952, 
         nx34954, nx34956, nx34958, nx34960, nx34962, nx34964, nx34966, nx34968, 
         nx34970, nx34972, nx34974, nx34976, nx34978, nx34980, nx34982, nx34984, 
         nx34986, nx34988, nx34990, nx34992, nx34994, nx34996, nx35004, nx35006, 
         nx35008, nx35010, nx35012, nx35014, nx35016, nx35018, nx35020, nx35022, 
         nx35024, nx35026, nx35028, nx35030, nx35032, nx35034, nx35036, nx35038, 
         nx35040, nx35042, nx35044, nx35046, nx35048, nx35050, nx35052, nx35054, 
         nx35056, nx35058, nx35060, nx35062, nx35064, nx35066, nx35074, nx35076, 
         nx35078, nx35080, nx35082, nx35084, nx35086, nx35088, nx35090, nx35092, 
         nx35094, nx35096, nx35098, nx35100, nx35102, nx35104, nx35106, nx35108, 
         nx35110, nx35112, nx35114, nx35116, nx35118, nx35120, nx35122, nx35124, 
         nx35126, nx35128, nx35130, nx35132, nx35134, nx35136, nx35140, nx35142, 
         nx35144, nx35146, nx35148, nx35150, nx35152, nx35154, nx35156, nx35158, 
         nx35160, nx35162, nx35164, nx35166, nx35168, nx35170, nx35172, nx35174, 
         nx35176, nx35178, nx35180, nx35182, nx35184, nx35186, nx35188, nx35190, 
         nx35192, nx35194, nx35196, nx35198, nx35200, nx35202, nx35204, nx35206, 
         nx35208, nx35210, nx35212, nx35216, nx35218, nx35220, nx35222, nx35224, 
         nx35226, nx35228, nx35230, nx35232, nx35234, nx35236, nx35238, nx35240, 
         nx35242, nx35244, nx35246, nx35248, nx35250, nx35252, nx35254, nx35256, 
         nx35258, nx35260, nx35262, nx35264, nx35266, nx35268, nx35270, nx35272, 
         nx35274, nx35276, nx35278, nx35280, nx35282, nx35284, nx35286, nx35288, 
         nx35292, nx35294, nx35296, nx35298, nx35300, nx35302, nx35304, nx35306, 
         nx35308, nx35310, nx35312, nx35314, nx35316, nx35318, nx35320, nx35322, 
         nx35324, nx35326, nx35328, nx35330, nx35332, nx35334, nx35336, nx35338, 
         nx35340, nx35342, nx35344, nx35346, nx35348, nx35350, nx35352, nx35354, 
         nx35356, nx35358, nx35360, nx35362, nx35364, nx35368, nx35370, nx35372, 
         nx35374, nx35376, nx35378, nx35380, nx35382, nx35384, nx35386, nx35388, 
         nx35390, nx35392, nx35394, nx35396, nx35398, nx35400, nx35402, nx35404, 
         nx35406, nx35408, nx35410, nx35412, nx35414, nx35416, nx35418, nx35420, 
         nx35422, nx35424, nx35426, nx35428, nx35430, nx35432, nx35434, nx35436, 
         nx35438, nx35440, nx35444, nx35446, nx35448, nx35450, nx35452, nx35454, 
         nx35456, nx35458, nx35460, nx35462, nx35464, nx35466, nx35468, nx35470, 
         nx35472, nx35474, nx35476, nx35478, nx35480, nx35482, nx35484, nx35486, 
         nx35488, nx35490, nx35492, nx35494, nx35496, nx35498, nx35500, nx35502, 
         nx35504, nx35506, nx35508, nx35510, nx35512, nx35514, nx35516, nx35520, 
         nx35522, nx35524, nx35526, nx35528, nx35530, nx35532, nx35534, nx35536, 
         nx35538, nx35540, nx35542, nx35544, nx35546, nx35548, nx35550, nx35552, 
         nx35554, nx35556, nx35558, nx35560, nx35562, nx35564, nx35566, nx35568, 
         nx35570, nx35572, nx35574, nx35576, nx35578, nx35580, nx35582, nx35584, 
         nx35586, nx35588, nx35590, nx35592, nx35596, nx35598, nx35600, nx35602, 
         nx35604, nx35606, nx35608, nx35610, nx35612, nx35614, nx35616, nx35618, 
         nx35620, nx35622, nx35624, nx35626, nx35628, nx35630, nx35632, nx35634, 
         nx35636, nx35638, nx35640, nx35642, nx35644, nx35646, nx35648, nx35650, 
         nx35652, nx35654, nx35656, nx35658, nx35660, nx35662, nx35664, nx35666, 
         nx35668, nx35670, nx35672, nx35674, nx35676, nx35678, nx35680, nx35682, 
         nx35684, nx35686, nx35688, nx35690, nx35692, nx35694, nx35696, nx35698, 
         nx35700, nx35702, nx35704, nx35706, nx35708, nx35712, nx35714, nx35716, 
         nx35718, nx35720, nx35782, nx35784, nx35786, nx35796, nx35798, nx35804, 
         nx35806, nx35808, nx35810, nx35812, nx35814, nx35816, nx35818, nx35820, 
         nx35822, nx35824, nx35826, nx35828, nx35830, nx35832, nx35834, nx35836, 
         nx35838, nx35840, nx35842, nx35844, nx35846, nx35848, nx35850, nx35852, 
         nx35854, nx35856, nx35858, nx35860, nx35862, nx35864, nx35866, nx35868, 
         nx35870, nx35872, nx35874, nx35876, nx35878, nx35880, nx35882, nx35884, 
         nx35886, nx35888, nx35890, nx35892, nx35894, nx35896, nx35898, nx35900, 
         nx35902, nx35904, nx35906, nx35908, nx35910, nx35912, nx35914, nx35916, 
         nx35918, nx35920, nx35922, nx35924, nx35926, nx35928, nx35930, nx35932, 
         nx35934, nx35936, nx35938, nx35940, nx35942, nx35944, nx35946, nx35948, 
         nx35950, nx35952, nx35954, nx35956, nx35958, nx35960, nx35962, nx35964, 
         nx35966, nx35968, nx35970, nx35972, nx35974, nx35976, nx35978, nx35980, 
         nx35982, nx35984, nx35986, nx35988, nx35990, nx35992, nx35994, nx35996, 
         nx35998, nx36000, nx36002, nx36004, nx36006, nx36008, nx36010, nx36012, 
         nx36014, nx36016, nx36018, nx36020, nx36022, nx36024, nx36026, nx36028, 
         nx36030, nx36032, nx36034, nx36036, nx36038, nx36040, nx36042, nx36044, 
         nx36046, nx36048, nx36050, nx36052, nx36054, nx36056, nx36058, nx36060, 
         nx36062, nx36064, nx36066, nx36068, nx36070, nx36072, nx36074, nx36076, 
         nx36078, nx36080, nx36082, nx36084, nx36086, nx36088, nx36090, nx36092, 
         nx36094, nx36096, nx36098, nx36100, nx36102, nx36104, nx36106, nx36108, 
         nx36110, nx36112, nx36114, nx36116, nx36118, nx36120, nx36122, nx36124, 
         nx36126, nx36128, nx36130, nx36132, nx36134, nx36136, nx36138, nx36140, 
         nx36142, nx36144, nx36146, nx36148, nx36150, nx36152, nx36154, nx36156, 
         nx36158, nx36160, nx36162, nx36164, nx36166, nx36168, nx36170, nx36172, 
         nx36174, nx36176, nx36178, nx36180, nx36182, nx36184, nx36186, nx36188, 
         nx36190, nx36192, nx36194, nx36196, nx36198, nx36200, nx36202, nx36204, 
         nx36206, nx36208, nx36210, nx36212, nx36214, nx36216, nx36218, nx36220, 
         nx36222, nx36224, nx36226, nx36228, nx36230, nx36232, nx36234, nx36236, 
         nx36238, nx36240, nx36242, nx36244, nx36246, nx36248, nx36250, nx36252, 
         nx36254, nx36256, nx36258, nx36260, nx36262, nx36264, nx36266, nx36268, 
         nx36270, nx36272, nx36274, nx36276, nx36278, nx36280, nx36282, nx36284, 
         nx36286, nx36288, nx36290, nx36292, nx36294, nx36296, nx36298, nx36300, 
         nx36302, nx36304, nx36306, nx36308, nx36310, nx36312, nx36314, nx36316, 
         nx36318, nx36320, nx36322, nx36324, nx36326, nx36328, nx36330, nx36332, 
         nx36334, nx36336, nx36338, nx36340, nx36342, nx36344, nx36346, nx36348, 
         nx36350, nx36352, nx36354, nx36356, nx36358, nx36360, nx36362, nx36364, 
         nx36366, nx36368, nx36370, nx36372, nx36374, nx36376, nx36378, nx36380, 
         nx36382, nx36384, nx36386, nx36388, nx36390, nx36392, nx36394, nx36396, 
         nx36398, nx36400, nx36402, nx36404, nx36406, nx36408, nx36410, nx36412, 
         nx36414, nx36416, nx36418, nx36420, nx36422, nx36424, nx36426, nx36428, 
         nx36430, nx36432, nx36434, nx36436, nx36438, nx36440, nx36442, nx36444, 
         nx36446, nx36448, nx36450, nx36452, nx36454, nx36456, nx36458, nx36460, 
         nx36462, nx36464, nx36466, nx36468, nx36470, nx36472, nx36474, nx36476, 
         nx36478, nx36480, nx36482, nx36484, nx36486, nx36488, nx36490, nx36492, 
         nx36494, nx36496, nx36498, nx36500, nx36506, nx36508, nx36510, nx36512, 
         nx36514, nx36516, nx36518, nx36520, nx36522, nx36524, nx36526, nx36528, 
         nx36530, nx36532, nx36534, nx36536, nx36538, nx36540, nx36542, nx36544, 
         nx36546, nx36548, nx36550, nx36552, nx36554, nx36556, nx36558, nx36560, 
         nx36562, nx36564, nx36566, nx36568, nx36570, nx36572, nx36574, nx36580, 
         nx36582, nx36584, nx36586, nx36588, nx36590, nx36592, nx36594, nx36596, 
         nx36598, nx36600, nx36602, nx36604, nx36606, nx36608, nx36610, nx36612, 
         nx36614, nx36616, nx36618, nx36620, nx36622, nx36624, nx36626, nx36628, 
         nx36630, nx36632, nx36634, nx36636, nx36638, nx36640, nx36642, nx36644, 
         nx36646, nx36648, nx36654, nx36656, nx36658, nx36660, nx36662, nx36664, 
         nx36666, nx36668, nx36670, nx36672, nx36674, nx36676, nx36678, nx36680, 
         nx36682, nx36684, nx36686, nx36688, nx36690, nx36692, nx36694, nx36696, 
         nx36698, nx36700, nx36702, nx36704, nx36706, nx36708, nx36710, nx36712, 
         nx36714, nx36716, nx36718, nx36720, nx36728, nx36730, nx36732, nx36734, 
         nx36736, nx36738, nx36740, nx36742, nx36744, nx36746, nx36748, nx36750, 
         nx36752, nx36754, nx36756, nx36758, nx36760, nx36762, nx36764, nx36766, 
         nx36768, nx36770, nx36772, nx36774, nx36776, nx36778, nx36780, nx36782, 
         nx36784, nx36786, nx36788, nx36790, nx36792, nx36794, nx36796, nx36804, 
         nx36806, nx36808, nx36810, nx36812, nx36814, nx36816, nx36818, nx36820, 
         nx36822, nx36824, nx36826, nx36828, nx36830, nx36832, nx36834, nx36836, 
         nx36838, nx36840, nx36842, nx36844, nx36846, nx36848, nx36850, nx36852, 
         nx36854, nx36856, nx36858, nx36860, nx36862, nx36864, nx36866, nx36868, 
         nx36870, nx36872, nx36874, nx36876, nx36878, nx36880, nx36882, nx36884, 
         nx36886, nx36888, nx36890, nx36892, nx36894, nx36896, nx36898, nx36912, 
         nx36916, nx36918, nx36920, nx36922, nx36924, nx36926, nx36928, nx36930, 
         nx36932, nx36934, nx36936, nx36938, nx36940, nx36942, nx36944, nx36946, 
         nx36948, nx36950, nx36952, nx36954, nx36956, nx36958, nx36960, nx36962, 
         nx36964, nx36966, nx36968, nx36970, nx36972, nx36974, nx36976, nx36978, 
         nx36980, nx36982, nx36984, nx36986, nx36988, nx36990, nx36992, nx36994, 
         nx36996, nx36998, nx37000, nx37002, nx37004, nx37006, nx37008, nx37010, 
         nx37012, nx37014, nx37016, nx37018, nx37020, nx37022, nx37024, nx37026, 
         nx37028, nx37030, nx37032, nx37034, nx37036, nx37038, nx37040, nx37042, 
         nx37044, nx37046, nx37048, nx37050, nx37052, nx37058, nx37060, nx37062, 
         nx37064, nx37066, nx37068, nx37070, nx37072, nx37074, nx37076, nx37078, 
         nx37080, nx37082, nx37084, nx37086, nx37088, nx37090, nx37092, nx37094, 
         nx37096, nx37098, nx37100, nx37102, nx37104, nx37106, nx37108, nx37110, 
         nx37112, nx37114, nx37116, nx37118, nx37120, nx37122, nx37124, nx37126, 
         nx37128, nx37130, nx37132, nx37134, nx37136, nx37138, nx37140, nx37142, 
         nx37144, nx37146, nx37148, nx37150, nx37152, nx37154, nx37156, nx37158, 
         nx37160, nx37162, nx37164, nx37166, nx37168, nx37170, nx37172, nx37174, 
         nx37176, nx37178, nx37180, nx37182, nx37184, nx37186, nx37188, nx37190, 
         nx37192, nx37194, nx37196, nx37198, nx37200, nx37202, nx37204, nx37206, 
         nx37208, nx37210, nx37212, nx37214, nx37216, nx37218, nx37220, nx37222, 
         nx37224, nx37226, nx37228, nx37230, nx37232, nx37234, nx37236, nx37238, 
         nx37240, nx37242, nx37244, nx37246, nx37248, nx37250, nx37252, nx37254, 
         nx37256, nx37258, nx37260, nx37262, nx37264, nx37266, nx37268, nx37270, 
         nx37272, nx37274, nx37276, nx37278, nx37280, nx37282, nx37284, nx37286, 
         nx37288, nx37290, nx37292, nx37294, nx37296, nx37298, nx37300, nx37302, 
         nx37304, nx37306, nx37308, nx37310, nx37312, nx37314, nx37316, nx37318, 
         nx37320, nx37322, nx37324, nx37326, nx37328, nx37330, nx37332, nx37334, 
         nx37336, nx37338, nx37340, nx37342, nx37344, nx37346, nx37348, nx37350, 
         nx37352, nx37354, nx37356, nx37358, nx37360, nx37362, nx37364, nx37366, 
         nx37368, nx37370, nx37372, nx37374, nx37376, nx37378, nx37380, nx37382, 
         nx37384, nx37386, nx37388, nx37390, nx37392, nx37394, nx37396, nx37398, 
         nx37400, nx37402, nx37404, nx37406, nx37412, nx37414, nx37416, nx37418, 
         nx37420, nx37422, nx37424, nx37426, nx37428, nx37430, nx37436, nx37438;
    wire [2112:0] \$dummy ;




    dff camera_module_algo_module_direc_reg_reg_q_0 (.Q (motor_direction[0]), .QB (
        \$dummy [0]), .D (nx22543), .CLK (clk)) ;
    mux21_ni ix22544 (.Y (nx22543), .A0 (motor_direction[0]), .A1 (nx27166), .S0 (
             nx27156)) ;
    oai21 ix1134 (.Y (nx1133), .A0 (nx35686), .A1 (nx34038), .B0 (nx34027)) ;
    dff camera_module_algo_module_modCU_reg_current_state_0 (.Q (
        camera_module_algo_module_regs_rst), .QB (\$dummy [1]), .D (nx1133), .CLK (
        clk)) ;
    nor03_2x ix1222 (.Y (nx1221), .A0 (nx22568), .A1 (rst), .A2 (nx33608)) ;
    nand03 ix22569 (.Y (nx22568), .A0 (nx512), .A1 (nx23021), .A2 (nx622)) ;
    nor03_2x ix513 (.Y (nx512), .A0 (camera_module_algo_module_address_value_1)
             , .A1 (camera_module_algo_module_address_value_3), .A2 (
             camera_module_algo_module_address_value_2)) ;
    mux21_ni ix1154 (.Y (nx1153), .A0 (nx448), .A1 (
             camera_module_algo_module_address_value_1), .S0 (nx22973)) ;
    oai32 ix449 (.Y (nx448), .A0 (nx22575), .A1 (nx34138), .A2 (
          camera_module_algo_module_prev_cont_enable), .B0 (nx35684), .B1 (
          nx35796)) ;
    xnor2 ix22576 (.Y (nx22575), .A0 (nx22577), .A1 (nx22931)) ;
    mux21_ni ix22578 (.Y (nx22577), .A0 (nx37094), .A1 (nx23021), .S0 (one)) ;
    oai21 ix1074 (.Y (nx1073), .A0 (nx22585), .A1 (nx34036), .B0 (nx22587)) ;
    dff camera_module_algo_module_modCU_reg_current_state_6 (.Q (
        camera_module_algo_module_modCU_current_state_6), .QB (nx22585), .D (
        nx1073), .CLK (clk)) ;
    oai22 ix1064 (.Y (nx1063), .A0 (nx22595), .A1 (nx34036), .B0 (rst), .B1 (
          nx22597)) ;
    dff camera_module_algo_module_modCU_reg_current_state_5 (.Q (
        camera_module_algo_module_modCU_current_state_5), .QB (nx22595), .D (
        nx1063), .CLK (clk)) ;
    oai22 ix1054 (.Y (nx1053), .A0 (nx22597), .A1 (nx34036), .B0 (rst), .B1 (
          nx22601)) ;
    nor02_2x ix309 (.Y (nx308), .A0 (rst), .A1 (nx22605)) ;
    aoi22 ix22606 (.Y (nx22605), .A0 (
          camera_module_algo_module_nvm_address_enable), .A1 (
          camera_module_ack_from_DMA), .B0 (
          camera_module_algo_module_modCU_current_state_12), .B1 (nx22568)) ;
    oai22 ix954 (.Y (nx953), .A0 (nx22611), .A1 (nx34036), .B0 (rst), .B1 (
          nx22613)) ;
    dff camera_module_algo_module_modCU_reg_current_state_2 (.Q (
        camera_module_algo_module_nvm_address_enable), .QB (nx22611), .D (nx953)
        , .CLK (clk)) ;
    aoi21 ix22614 (.Y (nx22613), .A0 (start), .A1 (
          camera_module_algo_module_modCU_current_state_1), .B0 (
          camera_module_algo_module_prev_cont_enable)) ;
    dff camera_module_algo_module_modCU_reg_current_state_1 (.Q (
        camera_module_algo_module_modCU_current_state_1), .QB (\$dummy [2]), .D (
        nx22523), .CLK (clk)) ;
    dff camera_module_algo_module_modCU_reg_current_state_13 (.Q (
        camera_module_algo_module_modCU_current_state_13), .QB (nx22565), .D (
        nx1221), .CLK (clk)) ;
    dff camera_module_algo_module_modCU_reg_current_state_14 (.Q (
        camera_module_algo_module_modCU_current_state_14), .QB (\$dummy [3]), .D (
        nx22481), .CLK (clk)) ;
    nor03_2x ix22482 (.Y (nx22481), .A0 (nx22627), .A1 (rst), .A2 (nx22565)) ;
    xnor2 ix22628 (.Y (nx22627), .A0 (nx26956), .A1 (nx27038)) ;
    oai22 ix26957 (.Y (nx26956), .A0 (nx22631), .A1 (nx33816), .B0 (nx33810), .B1 (
          camera_module_algo_module_prev_cont_value_15)) ;
    dff camera_module_algo_module_curr_cont_reg_reg_q_15 (.Q (
        camera_module_algo_module_current_cont_value_15), .QB (nx33810), .D (
        nx22273), .CLK (clk)) ;
    dff camera_module_algo_module_Addout_reg_reg_q_15 (.Q (
        camera_module_algo_module_Addout_value_15), .QB (\$dummy [4]), .D (
        nx22263), .CLK (clk)) ;
    xnor2 ix26545 (.Y (nx26544), .A0 (nx26504), .A1 (nx33790)) ;
    oai22 ix26505 (.Y (nx26504), .A0 (nx22645), .A1 (nx33765), .B0 (nx33779), .B1 (
          nx33776)) ;
    aoi22 ix22646 (.Y (nx22645), .A0 (camera_module_algo_module_diff_value_13), 
          .A1 (camera_module_algo_module_current_cont_value_13), .B0 (nx26356), 
          .B1 (nx933)) ;
    dff camera_module_algo_module_diff_reg_reg_q_13 (.Q (
        camera_module_algo_module_diff_value_13), .QB (nx22651), .D (nx22213), .CLK (
        clk)) ;
    aoi21 ix22654 (.Y (nx22653), .A0 (zero), .A1 (nx34118), .B0 (nx26412)) ;
    nor03_2x ix26413 (.Y (nx26412), .A0 (nx34118), .A1 (nx35700), .A2 (nx33384)
             ) ;
    mux21_ni ix1254 (.Y (nx1253), .A0 (zero), .A1 (
             camera_module_algo_module_pixel_value_8), .S0 (nx37152)) ;
    dff camera_module_algo_module_pixel_reg_reg_q_8 (.Q (
        camera_module_algo_module_pixel_value_8), .QB (\$dummy [5]), .D (nx1253)
        , .CLK (clk)) ;
    dff camera_module_algo_module_modCU_reg_current_state_3 (.Q (
        camera_module_algo_module_pixel_enable), .QB (nx22601), .D (nx1043), .CLK (
        clk)) ;
    aoi21 ix22670 (.Y (nx22669), .A0 (nx37086), .A1 (nx25422), .B0 (nx704)) ;
    oai21 ix25423 (.Y (nx25422), .A0 (nx35708), .A1 (nx22681), .B0 (nx22679)) ;
    oai21 ix22678 (.Y (nx22677), .A0 (camera_module_algo_module_pixel_value_8), 
          .A1 (nx35670), .B0 (nx22679)) ;
    nand02 ix22680 (.Y (nx22679), .A0 (nx35670), .A1 (
           camera_module_algo_module_pixel_value_8)) ;
    aoi21 ix22682 (.Y (nx22681), .A0 (nx37086), .A1 (nx25414), .B0 (nx704)) ;
    oai21 ix25415 (.Y (nx25414), .A0 (nx35708), .A1 (nx22685), .B0 (nx22679)) ;
    aoi21 ix22686 (.Y (nx22685), .A0 (nx37086), .A1 (nx25406), .B0 (nx704)) ;
    oai21 ix25407 (.Y (nx25406), .A0 (nx35708), .A1 (nx22689), .B0 (nx22679)) ;
    aoi21 ix22690 (.Y (nx22689), .A0 (nx25398), .A1 (nx37086), .B0 (nx704)) ;
    oai22 ix25399 (.Y (nx25398), .A0 (nx22693), .A1 (nx32243), .B0 (nx33382), .B1 (
          nx25374)) ;
    aoi22 ix22694 (.Y (nx22693), .A0 (camera_module_algo_module_pixel_value_6), 
          .A1 (nx22699), .B0 (nx19850), .B1 (nx22616)) ;
    dff camera_module_algo_module_pixel_reg_reg_q_6 (.Q (
        camera_module_algo_module_pixel_value_6), .QB (\$dummy [6]), .D (nx19243
        ), .CLK (clk)) ;
    mux21_ni ix19244 (.Y (nx19243), .A0 (nx22608), .A1 (
             camera_module_algo_module_pixel_value_6), .S0 (nx37152)) ;
    mux21_ni ix22700 (.Y (nx22699), .A0 (nx22701), .A1 (nx35674), .S0 (nx36792)
             ) ;
    nor04 ix22702 (.Y (nx22701), .A0 (nx22588), .A1 (nx21934), .A2 (nx21278), .A3 (
          nx20624)) ;
    nand04 ix22589 (.Y (nx22588), .A0 (nx22705), .A1 (nx23302), .A2 (nx23413), .A3 (
           nx23520)) ;
    oai21 ix22706 (.Y (nx22705), .A0 (nx22578), .A1 (nx22500), .B0 (nx36448)) ;
    nand04 ix22579 (.Y (nx22578), .A0 (nx22709), .A1 (nx23138), .A2 (nx23165), .A3 (
           nx23189)) ;
    aoi22 ix22710 (.Y (nx22709), .A0 (camera_module_cache_ram_0__6), .A1 (
          nx37030), .B0 (camera_module_cache_ram_16__6), .B1 (nx37032)) ;
    dffr camera_module_cache_reg_ram_0__6 (.Q (camera_module_cache_ram_0__6), .QB (
         \$dummy [7]), .D (nx19233), .CLK (clk), .R (rst)) ;
    mux21_ni ix19234 (.Y (nx19233), .A0 (camera_module_cache_ram_0__6), .A1 (
             nx35520), .S0 (nx35134)) ;
    oai221 ix19971 (.Y (nx19970), .A0 (nx34072), .A1 (nx22851), .B0 (nx22871), .B1 (
           nx35712), .C0 (nx22874)) ;
    oai32 ix994 (.Y (nx993), .A0 (nx22719), .A1 (nx34070), .A2 (nx34042), .B0 (
          nx22846), .B1 (nx22779)) ;
    dff camera_module_DMA_module_R_Cache_addr_reg_q_3 (.Q (\$dummy [8]), .QB (
        nx22719), .D (nx993), .CLK (clk)) ;
    dff camera_module_DMA_module_controlUnit_reg_state_0 (.Q (
        camera_module_DMA_module_signals_1), .QB (\$dummy [9]), .D (nx20), .CLK (
        clk)) ;
    dff camera_module_DMA_module_controlUnit_reg_state_5 (.Q (
        camera_module_ack_from_DMA), .QB (nx22844), .D (nx294), .CLK (clk)) ;
    nor03_2x ix295 (.Y (nx294), .A0 (nx22727), .A1 (rst), .A2 (nx22795)) ;
    nand04 ix22728 (.Y (nx22727), .A0 (camera_module_cache_address_from_DMA_7), 
           .A1 (camera_module_cache_address_from_DMA_6), .A2 (
           camera_module_cache_address_from_DMA_5), .A3 (
           camera_module_cache_address_from_DMA_4)) ;
    dff camera_module_DMA_module_R_Cache_addr_reg_q_7 (.Q (
        camera_module_cache_address_from_DMA_7), .QB (\$dummy [10]), .D (nx1033)
        , .CLK (clk)) ;
    mux21_ni ix1034 (.Y (nx1033), .A0 (nx276), .A1 (
             camera_module_cache_address_from_DMA_7), .S0 (nx22779)) ;
    xnor2 ix269 (.Y (nx268), .A0 (nx264), .A1 (nx22841)) ;
    oai22 ix265 (.Y (nx264), .A0 (nx22739), .A1 (nx22831), .B0 (nx35672), .B1 (
          nx22835)) ;
    aoi22 ix22740 (.Y (nx22739), .A0 (zero), .A1 (
          camera_module_cache_address_from_DMA_5), .B0 (nx216), .B1 (nx897)) ;
    dff camera_module_DMA_module_R_Cache_addr_reg_q_5 (.Q (
        camera_module_cache_address_from_DMA_5), .QB (\$dummy [11]), .D (nx1013)
        , .CLK (clk)) ;
    mux21_ni ix1014 (.Y (nx1013), .A0 (nx226), .A1 (
             camera_module_cache_address_from_DMA_5), .S0 (nx37154)) ;
    xnor2 ix219 (.Y (nx218), .A0 (nx216), .A1 (nx22827)) ;
    oai22 ix217 (.Y (nx216), .A0 (nx22749), .A1 (nx22815), .B0 (nx35672), .B1 (
          nx22821)) ;
    aoi22 ix22750 (.Y (nx22749), .A0 (zero), .A1 (nx34072), .B0 (nx126), .B1 (
          nx128)) ;
    oai22 ix127 (.Y (nx126), .A0 (nx22753), .A1 (nx22777), .B0 (nx35670), .B1 (
          nx37106)) ;
    aoi22 ix22754 (.Y (nx22753), .A0 (zero), .A1 (nx34098), .B0 (nx78), .B1 (
          nx889)) ;
    oai32 ix974 (.Y (nx973), .A0 (nx37096), .A1 (nx34066), .A2 (nx34040), .B0 (
          nx22805), .B1 (nx37154)) ;
    dff camera_module_DMA_module_R_Cache_addr_reg_q_1 (.Q (\$dummy [12]), .QB (
        nx22757), .D (nx973), .CLK (clk)) ;
    nor02_2x ix179 (.Y (nx178), .A0 (rst), .A1 (nx22761)) ;
    aoi221 ix22762 (.Y (nx22761), .A0 (
           camera_module_DMA_module_controlUnit_state_4), .A1 (nx22727), .B0 (
           nx34040), .B1 (nx35712), .C0 (camera_module_DMA_module_signals_4)) ;
    dff camera_module_DMA_module_controlUnit_reg_state_4 (.Q (
        camera_module_DMA_module_controlUnit_state_4), .QB (nx22795), .D (nx160)
        , .CLK (clk)) ;
    nor03_2x ix161 (.Y (nx160), .A0 (nx35712), .A1 (rst), .A2 (nx37028)) ;
    oai32 ix984 (.Y (nx983), .A0 (nx37106), .A1 (nx34066), .A2 (nx34040), .B0 (
          nx22773), .B1 (nx37154)) ;
    dff camera_module_DMA_module_R_Cache_addr_reg_q_2 (.Q (\$dummy [13]), .QB (
        nx22771), .D (nx983), .CLK (clk)) ;
    xnor2 ix22776 (.Y (nx22775), .A0 (nx22753), .A1 (nx22777)) ;
    oai32 ix964 (.Y (nx963), .A0 (nx37156), .A1 (nx34066), .A2 (nx34040), .B0 (
          nx22787), .B1 (nx37154)) ;
    dff camera_module_DMA_module_R_Cache_addr_reg_q_0 (.Q (
        camera_module_cache_address_from_DMA_0), .QB (\$dummy [14]), .D (nx963)
        , .CLK (clk)) ;
    xnor2 ix57 (.Y (nx56), .A0 (one), .A1 (nx22791)) ;
    dff camera_module_DMA_module_controlUnit_reg_state_3 (.Q (
        camera_module_write_from_DMA), .QB (\$dummy [15]), .D (nx178), .CLK (clk
        )) ;
    dff camera_module_DMA_module_controlUnit_reg_state_2 (.Q (
        camera_module_DMA_module_signals_4), .QB (\$dummy [16]), .D (nx48), .CLK (
        clk)) ;
    dff camera_module_DMA_module_controlUnit_reg_state_1 (.Q (
        camera_module_DMA_module_controlUnit_state_1), .QB (\$dummy [17]), .D (
        nx36), .CLK (clk)) ;
    nor02_2x ix37 (.Y (nx36), .A0 (rst), .A1 (nx22801)) ;
    aoi21 ix22802 (.Y (nx22801), .A0 (nx22611), .A1 (
          camera_module_DMA_module_controlUnit_state_1), .B0 (nx34066)) ;
    xnor2 ix81 (.Y (nx80), .A0 (nx78), .A1 (nx22811)) ;
    oai32 ix1004 (.Y (nx1003), .A0 (nx22821), .A1 (nx34068), .A2 (nx34040), .B0 (
          nx22823), .B1 (nx37154)) ;
    dff camera_module_DMA_module_R_Cache_addr_reg_q_4 (.Q (
        camera_module_cache_address_from_DMA_4), .QB (nx22821), .D (nx1003), .CLK (
        clk)) ;
    xnor2 ix22826 (.Y (nx22825), .A0 (nx22749), .A1 (nx22815)) ;
    xnor2 ix22828 (.Y (nx22827), .A0 (camera_module_cache_address_from_DMA_5), .A1 (
          zero)) ;
    oai32 ix1024 (.Y (nx1023), .A0 (nx22835), .A1 (nx34068), .A2 (nx34040), .B0 (
          nx22837), .B1 (nx37154)) ;
    dff camera_module_DMA_module_R_Cache_addr_reg_q_6 (.Q (
        camera_module_cache_address_from_DMA_6), .QB (nx22835), .D (nx1023), .CLK (
        clk)) ;
    xnor2 ix22840 (.Y (nx22839), .A0 (nx22739), .A1 (nx22831)) ;
    xnor2 ix22842 (.Y (nx22841), .A0 (camera_module_cache_address_from_DMA_7), .A1 (
          zero)) ;
    xnor2 ix131 (.Y (nx130), .A0 (nx126), .A1 (nx22849)) ;
    tri01 nvm_module_tri_dataout_126 (.Y (nvm_data_126), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_118 (.Y (nvm_data_118), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_110 (.Y (nvm_data_110), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_102 (.Y (nvm_data_102), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_94 (.Y (nvm_data_94), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_86 (.Y (nvm_data_86), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_78 (.Y (nvm_data_78), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_70 (.Y (nvm_data_70), .A (nx22549), .E (
          nvm_module_GND0)) ;
    inv01 ix22872 (.Y (nx22871), .A (nvm_data_6)) ;
    tri01 nvm_module_tri_dataout_6 (.Y (nvm_data_6), .A (nx22549), .E (
          nvm_module_GND0)) ;
    nand02 ix22875 (.Y (nx22874), .A0 (nx34072), .A1 (nx19904)) ;
    tri01 nvm_module_tri_dataout_62 (.Y (nvm_data_62), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_54 (.Y (nvm_data_54), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_46 (.Y (nvm_data_46), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_38 (.Y (nvm_data_38), .A (nx22549), .E (
          nvm_module_GND0)) ;
    oai22 ix19873 (.Y (nx19872), .A0 (nx34098), .A1 (nx22887), .B0 (nx34080), .B1 (
          nx22891)) ;
    tri01 nvm_module_tri_dataout_30 (.Y (nvm_data_30), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_22 (.Y (nvm_data_22), .A (nx22549), .E (
          nvm_module_GND0)) ;
    nand02 ix22892 (.Y (nx22891), .A0 (nvm_data_14), .A1 (nx34100)) ;
    tri01 nvm_module_tri_dataout_14 (.Y (nvm_data_14), .A (nx22549), .E (
          nvm_module_GND0)) ;
    nand02 ix1491 (.Y (nx1490), .A0 (nx22897), .A1 (nx23073)) ;
    nor02_2x ix22898 (.Y (nx22897), .A0 (nx1050), .A1 (nx1024)) ;
    xnor2 ix1039 (.Y (nx1038), .A0 (nx1004), .A1 (nx23033)) ;
    oai22 ix1005 (.Y (nx1004), .A0 (nx22907), .A1 (nx23012), .B0 (nx23011), .B1 (
          nx37196)) ;
    dff camera_module_algo_module_Address_reg_reg_q_5 (.Q (
        camera_module_algo_module_address_value_5), .QB (nx23011), .D (nx1193), 
        .CLK (clk)) ;
    mux21_ni ix1194 (.Y (nx1193), .A0 (nx552), .A1 (
             camera_module_algo_module_address_value_5), .S0 (nx37198)) ;
    oai32 ix553 (.Y (nx552), .A0 (nx22912), .A1 (nx34120), .A2 (
          camera_module_algo_module_prev_cont_enable), .B0 (nx35672), .B1 (
          nx35786)) ;
    xnor2 ix22913 (.Y (nx22912), .A0 (nx22915), .A1 (nx22907)) ;
    aoi22 ix22916 (.Y (nx22915), .A0 (camera_module_algo_module_address_value_4)
          , .A1 (nx34140), .B0 (nx518), .B1 (nx905)) ;
    dff camera_module_algo_module_Address_reg_reg_q_4 (.Q (
        camera_module_algo_module_address_value_4), .QB (\$dummy [18]), .D (
        nx1183), .CLK (clk)) ;
    mux21_ni ix1184 (.Y (nx1183), .A0 (nx528), .A1 (
             camera_module_algo_module_address_value_4), .S0 (nx37198)) ;
    xnor2 ix521 (.Y (nx520), .A0 (nx518), .A1 (nx23006)) ;
    oai22 ix519 (.Y (nx518), .A0 (nx22923), .A1 (nx22997), .B0 (nx23005), .B1 (
          nx37196)) ;
    aoi22 ix22924 (.Y (nx22923), .A0 (camera_module_algo_module_address_value_2)
          , .A1 (nx34140), .B0 (nx460), .B1 (nx903)) ;
    dff camera_module_algo_module_Address_reg_reg_q_2 (.Q (
        camera_module_algo_module_address_value_2), .QB (\$dummy [19]), .D (
        nx1163), .CLK (clk)) ;
    mux21_ni ix1164 (.Y (nx1163), .A0 (nx470), .A1 (
             camera_module_algo_module_address_value_2), .S0 (nx37198)) ;
    xnor2 ix463 (.Y (nx462), .A0 (nx460), .A1 (nx22951)) ;
    oai22 ix461 (.Y (nx460), .A0 (nx22577), .A1 (nx22931), .B0 (nx22935), .B1 (
          nx37196)) ;
    xnor2 ix437 (.Y (nx436), .A0 (zero), .A1 (nx37094)) ;
    dff camera_module_algo_module_Address_reg_reg_q_1 (.Q (
        camera_module_algo_module_address_value_1), .QB (nx22935), .D (nx1153), 
        .CLK (clk)) ;
    oai21 ix1094 (.Y (nx1093), .A0 (nx22943), .A1 (nx34036), .B0 (nx22945)) ;
    dff camera_module_algo_module_modCU_reg_current_state_8 (.Q (\$dummy [20]), 
        .QB (nx22943), .D (nx1093), .CLK (clk)) ;
    nand03 ix22946 (.Y (nx22945), .A0 (nx35692), .A1 (
           camera_module_algo_module_modCU_current_state_7), .A2 (nx34036)) ;
    dff camera_module_algo_module_modCU_reg_current_state_7 (.Q (
        camera_module_algo_module_modCU_current_state_7), .QB (\$dummy [21]), .D (
        nx1083), .CLK (clk)) ;
    dff camera_module_algo_module_modCU_reg_current_state_16 (.Q (
        camera_module_algo_module_prev_cont_enable), .QB (\$dummy [22]), .D (
        nx22513), .CLK (clk)) ;
    ao32 ix22514 (.Y (nx22513), .A0 (motor_move), .A1 (motor_done), .A2 (nx35692
         ), .B0 (camera_module_algo_module_prev_cont_enable), .B1 (nx35696)) ;
    dff camera_module_algo_module_modCU_reg_current_state_15 (.Q (motor_move), .QB (
        \$dummy [23]), .D (nx22503), .CLK (clk)) ;
    nor02_2x ix27085 (.Y (nx27084), .A0 (rst), .A1 (nx22961)) ;
    aoi22 ix22962 (.Y (nx22961), .A0 (nx22963), .A1 (
          camera_module_algo_module_modCU_current_state_14), .B0 (
          camera_module_algo_module_modCU_current_state_13), .B1 (nx22627)) ;
    mux21_ni ix22494 (.Y (nx22493), .A0 (nx27068), .A1 (
             camera_module_algo_module_failure_count_value_0), .S0 (nx22968)) ;
    dff camera_module_algo_module_fail_count_reg_reg_q_0 (.Q (
        camera_module_algo_module_failure_count_value_0), .QB (nx22963), .D (
        nx22493), .CLK (clk)) ;
    nor03_2x ix22969 (.Y (nx22968), .A0 (
             camera_module_algo_module_modCU_current_state_14), .A1 (motor_move)
             , .A2 (nx34118)) ;
    oai21 ix1124 (.Y (nx1123), .A0 (nx22979), .A1 (nx34036), .B0 (nx22981)) ;
    dff camera_module_algo_module_modCU_reg_current_state_11 (.Q (\$dummy [24])
        , .QB (nx22979), .D (nx1123), .CLK (clk)) ;
    oai21 ix1114 (.Y (nx1113), .A0 (nx22987), .A1 (nx34038), .B0 (nx22989)) ;
    dff camera_module_algo_module_modCU_reg_current_state_10 (.Q (
        camera_module_algo_module_modCU_current_state_10), .QB (nx22987), .D (
        nx1113), .CLK (clk)) ;
    oai22 ix1104 (.Y (nx1103), .A0 (nx22993), .A1 (nx34038), .B0 (rst), .B1 (
          nx22943)) ;
    dff camera_module_algo_module_modCU_reg_current_state_9 (.Q (\$dummy [25]), 
        .QB (nx22993), .D (nx1103), .CLK (clk)) ;
    dff camera_module_algo_module_Address_reg_reg_q_3 (.Q (
        camera_module_algo_module_address_value_3), .QB (nx23005), .D (nx1173), 
        .CLK (clk)) ;
    mux21_ni ix1174 (.Y (nx1173), .A0 (nx496), .A1 (
             camera_module_algo_module_address_value_3), .S0 (nx37198)) ;
    oai32 ix497 (.Y (nx496), .A0 (nx23003), .A1 (nx34118), .A2 (
          camera_module_algo_module_prev_cont_enable), .B0 (nx35672), .B1 (
          nx35786)) ;
    xnor2 ix23004 (.Y (nx23003), .A0 (nx22923), .A1 (nx22997)) ;
    aoi22 ix23013 (.Y (nx23012), .A0 (camera_module_algo_module_address_value_4)
          , .A1 (nx426), .B0 (nx932), .B1 (nx934)) ;
    xnor2 ix427 (.Y (nx426), .A0 (one), .A1 (nx37094)) ;
    oai22 ix933 (.Y (nx932), .A0 (nx22997), .A1 (nx23016), .B0 (nx23005), .B1 (
          nx37196)) ;
    aoi22 ix23017 (.Y (nx23016), .A0 (camera_module_algo_module_address_value_2)
          , .A1 (nx34142), .B0 (nx903), .B1 (nx860)) ;
    oai22 ix861 (.Y (nx860), .A0 (nx22935), .A1 (nx37196), .B0 (nx22931), .B1 (
          nx23019)) ;
    mux21_ni ix23020 (.Y (nx23019), .A0 (nx37094), .A1 (nx23021), .S0 (zero)) ;
    mux21_ni ix1144 (.Y (nx1143), .A0 (nx418), .A1 (
             camera_module_algo_module_address_value_0), .S0 (nx37198)) ;
    oai32 ix419 (.Y (nx418), .A0 (nx23026), .A1 (nx34120), .A2 (
          camera_module_algo_module_prev_cont_enable), .B0 (nx35672), .B1 (
          nx35786)) ;
    dff camera_module_algo_module_Address_reg_reg_q_0 (.Q (
        camera_module_algo_module_address_value_0), .QB (nx23021), .D (nx1143), 
        .CLK (clk)) ;
    dff camera_module_algo_module_Address_reg_reg_q_6 (.Q (
        camera_module_algo_module_address_value_6), .QB (\$dummy [26]), .D (
        nx1203), .CLK (clk)) ;
    mux21_ni ix1204 (.Y (nx1203), .A0 (nx576), .A1 (
             camera_module_algo_module_address_value_6), .S0 (nx37198)) ;
    xnor2 ix569 (.Y (nx568), .A0 (nx566), .A1 (nx23033)) ;
    oai22 ix567 (.Y (nx566), .A0 (nx22915), .A1 (nx22907), .B0 (nx23011), .B1 (
          nx37196)) ;
    dff camera_module_algo_module_modCU_reg_current_state_4 (.Q (\$dummy [27]), 
        .QB (nx22597), .D (nx1053), .CLK (clk)) ;
    oai32 ix1017 (.Y (nx1016), .A0 (
          camera_module_algo_module_modCU_current_state_6), .A1 (
          camera_module_algo_module_modCU_current_state_10), .A2 (nx23051), .B0 (
          nx35804), .B1 (nx23069)) ;
    xnor2 ix23054 (.Y (nx23053), .A0 (nx23055), .A1 (nx23059)) ;
    aoi22 ix23056 (.Y (nx23055), .A0 (camera_module_algo_module_address_value_6)
          , .A1 (nx34142), .B0 (nx566), .B1 (nx908)) ;
    dff camera_module_algo_module_Address_reg_reg_q_7 (.Q (
        camera_module_algo_module_address_value_7), .QB (nx23067), .D (nx1213), 
        .CLK (clk)) ;
    mux21_ni ix1214 (.Y (nx1213), .A0 (nx602), .A1 (
             camera_module_algo_module_address_value_7), .S0 (nx22973)) ;
    oai32 ix603 (.Y (nx602), .A0 (nx23053), .A1 (nx34120), .A2 (
          camera_module_algo_module_prev_cont_enable), .B0 (nx35672), .B1 (
          nx35786)) ;
    xnor2 ix23070 (.Y (nx23069), .A0 (nx23071), .A1 (nx23059)) ;
    aoi22 ix23072 (.Y (nx23071), .A0 (camera_module_algo_module_address_value_6)
          , .A1 (nx34142), .B0 (nx908), .B1 (nx1004)) ;
    nor02_2x ix23074 (.Y (nx23073), .A0 (nx980), .A1 (nx954)) ;
    xnor2 ix969 (.Y (nx968), .A0 (nx932), .A1 (nx23079)) ;
    xnor2 ix23080 (.Y (nx23079), .A0 (camera_module_algo_module_address_value_4)
          , .A1 (nx426)) ;
    oai32 ix947 (.Y (nx946), .A0 (
          camera_module_algo_module_modCU_current_state_6), .A1 (
          camera_module_algo_module_modCU_current_state_10), .A2 (nx23084), .B0 (
          nx35804), .B1 (nx23087)) ;
    xnor2 ix23088 (.Y (nx23087), .A0 (nx23012), .A1 (nx22907)) ;
    nand02 ix5651 (.Y (nx5650), .A0 (nx23091), .A1 (nx23105)) ;
    nor02_2x ix23092 (.Y (nx23091), .A0 (nx906), .A1 (nx880)) ;
    xnor2 ix895 (.Y (nx894), .A0 (nx860), .A1 (nx22951)) ;
    oai32 ix873 (.Y (nx872), .A0 (
          camera_module_algo_module_modCU_current_state_6), .A1 (
          camera_module_algo_module_modCU_current_state_10), .A2 (nx23100), .B0 (
          nx35804), .B1 (nx23102)) ;
    xnor2 ix23103 (.Y (nx23102), .A0 (nx23016), .A1 (nx22997)) ;
    nor02_2x ix23106 (.Y (nx23105), .A0 (nx836), .A1 (nx810)) ;
    oai32 ix829 (.Y (nx828), .A0 (
          camera_module_algo_module_modCU_current_state_6), .A1 (
          camera_module_algo_module_modCU_current_state_10), .A2 (nx23111), .B0 (
          nx35804), .B1 (nx23113)) ;
    oai32 ix803 (.Y (nx802), .A0 (
          camera_module_algo_module_modCU_current_state_6), .A1 (
          camera_module_algo_module_modCU_current_state_10), .A2 (nx23117), .B0 (
          nx23119), .B1 (nx35806)) ;
    xnor2 ix23120 (.Y (nx23119), .A0 (nx23019), .A1 (nx22931)) ;
    dffr camera_module_cache_reg_ram_16__6 (.Q (camera_module_cache_ram_16__6), 
         .QB (\$dummy [28]), .D (nx19223), .CLK (clk), .R (rst)) ;
    mux21_ni ix19224 (.Y (nx19223), .A0 (camera_module_cache_ram_16__6), .A1 (
             nx35520), .S0 (nx35130)) ;
    nand02 ix1473 (.Y (nx1472), .A0 (nx23130), .A1 (nx22897)) ;
    aoi22 ix23139 (.Y (nx23138), .A0 (camera_module_cache_ram_32__6), .A1 (
          nx37034), .B0 (camera_module_cache_ram_48__6), .B1 (nx37036)) ;
    dffr camera_module_cache_reg_ram_32__6 (.Q (camera_module_cache_ram_32__6), 
         .QB (\$dummy [29]), .D (nx19213), .CLK (clk), .R (rst)) ;
    mux21_ni ix19214 (.Y (nx19213), .A0 (camera_module_cache_ram_32__6), .A1 (
             nx35520), .S0 (nx35126)) ;
    nand02 ix1453 (.Y (nx1452), .A0 (nx23145), .A1 (nx22897)) ;
    dffr camera_module_cache_reg_ram_48__6 (.Q (camera_module_cache_ram_48__6), 
         .QB (\$dummy [30]), .D (nx19203), .CLK (clk), .R (rst)) ;
    mux21_ni ix19204 (.Y (nx19203), .A0 (camera_module_cache_ram_48__6), .A1 (
             nx35520), .S0 (nx35122)) ;
    nand02 ix1435 (.Y (nx1434), .A0 (nx23157), .A1 (nx22897)) ;
    nand02 ix987 (.Y (nx986), .A0 (nx980), .A1 (nx954)) ;
    aoi22 ix23166 (.Y (nx23165), .A0 (camera_module_cache_ram_64__6), .A1 (
          nx37038), .B0 (camera_module_cache_ram_80__6), .B1 (nx37040)) ;
    dffr camera_module_cache_reg_ram_64__6 (.Q (camera_module_cache_ram_64__6), 
         .QB (\$dummy [31]), .D (nx19193), .CLK (clk), .R (rst)) ;
    mux21_ni ix19194 (.Y (nx19193), .A0 (camera_module_cache_ram_64__6), .A1 (
             nx35520), .S0 (nx35118)) ;
    nand02 ix1411 (.Y (nx1410), .A0 (nx23172), .A1 (nx23073)) ;
    dffr camera_module_cache_reg_ram_80__6 (.Q (camera_module_cache_ram_80__6), 
         .QB (\$dummy [32]), .D (nx19183), .CLK (clk), .R (rst)) ;
    mux21_ni ix19184 (.Y (nx19183), .A0 (camera_module_cache_ram_80__6), .A1 (
             nx35520), .S0 (nx35114)) ;
    nand02 ix1393 (.Y (nx1392), .A0 (nx23172), .A1 (nx23130)) ;
    aoi22 ix23190 (.Y (nx23189), .A0 (camera_module_cache_ram_112__6), .A1 (
          nx37042), .B0 (camera_module_cache_ram_96__6), .B1 (nx37044)) ;
    dffr camera_module_cache_reg_ram_112__6 (.Q (camera_module_cache_ram_112__6)
         , .QB (\$dummy [33]), .D (nx19163), .CLK (clk), .R (rst)) ;
    mux21_ni ix19164 (.Y (nx19163), .A0 (camera_module_cache_ram_112__6), .A1 (
             nx35520), .S0 (nx35106)) ;
    nand02 ix1355 (.Y (nx1354), .A0 (nx23172), .A1 (nx23157)) ;
    dffr camera_module_cache_reg_ram_96__6 (.Q (camera_module_cache_ram_96__6), 
         .QB (\$dummy [34]), .D (nx19173), .CLK (clk), .R (rst)) ;
    mux21_ni ix19174 (.Y (nx19173), .A0 (camera_module_cache_ram_96__6), .A1 (
             nx35522), .S0 (nx35110)) ;
    nand02 ix1373 (.Y (nx1372), .A0 (nx23172), .A1 (nx23145)) ;
    nand04 ix22501 (.Y (nx22500), .A0 (nx23211), .A1 (nx23236), .A2 (nx23256), .A3 (
           nx23282)) ;
    aoi22 ix23212 (.Y (nx23211), .A0 (camera_module_cache_ram_128__6), .A1 (
          nx37046), .B0 (camera_module_cache_ram_144__6), .B1 (nx37048)) ;
    dffr camera_module_cache_reg_ram_128__6 (.Q (camera_module_cache_ram_128__6)
         , .QB (\$dummy [35]), .D (nx19153), .CLK (clk), .R (rst)) ;
    mux21_ni ix19154 (.Y (nx19153), .A0 (camera_module_cache_ram_128__6), .A1 (
             nx35522), .S0 (nx35102)) ;
    nand02 ix1327 (.Y (nx1326), .A0 (nx23218), .A1 (nx23073)) ;
    dffr camera_module_cache_reg_ram_144__6 (.Q (camera_module_cache_ram_144__6)
         , .QB (\$dummy [36]), .D (nx19143), .CLK (clk), .R (rst)) ;
    mux21_ni ix19144 (.Y (nx19143), .A0 (camera_module_cache_ram_144__6), .A1 (
             nx35522), .S0 (nx35098)) ;
    nand02 ix1309 (.Y (nx1308), .A0 (nx23218), .A1 (nx23130)) ;
    aoi22 ix23237 (.Y (nx23236), .A0 (camera_module_cache_ram_176__6), .A1 (
          nx37050), .B0 (camera_module_cache_ram_160__6), .B1 (nx37052)) ;
    dffr camera_module_cache_reg_ram_176__6 (.Q (camera_module_cache_ram_176__6)
         , .QB (\$dummy [37]), .D (nx19123), .CLK (clk), .R (rst)) ;
    mux21_ni ix19124 (.Y (nx19123), .A0 (camera_module_cache_ram_176__6), .A1 (
             nx35522), .S0 (nx35090)) ;
    nand02 ix1271 (.Y (nx1270), .A0 (nx23218), .A1 (nx23157)) ;
    dffr camera_module_cache_reg_ram_160__6 (.Q (camera_module_cache_ram_160__6)
         , .QB (\$dummy [38]), .D (nx19133), .CLK (clk), .R (rst)) ;
    mux21_ni ix19134 (.Y (nx19133), .A0 (camera_module_cache_ram_160__6), .A1 (
             nx35522), .S0 (nx35094)) ;
    nand02 ix1289 (.Y (nx1288), .A0 (nx23218), .A1 (nx23145)) ;
    aoi22 ix23257 (.Y (nx23256), .A0 (camera_module_cache_ram_192__6), .A1 (
          nx36288), .B0 (camera_module_cache_ram_208__6), .B1 (nx36328)) ;
    dffr camera_module_cache_reg_ram_192__6 (.Q (camera_module_cache_ram_192__6)
         , .QB (\$dummy [39]), .D (nx19113), .CLK (clk), .R (rst)) ;
    mux21_ni ix19114 (.Y (nx19113), .A0 (camera_module_cache_ram_192__6), .A1 (
             nx35522), .S0 (nx35086)) ;
    nand02 ix1057 (.Y (nx1056), .A0 (nx1050), .A1 (nx1024)) ;
    dffr camera_module_cache_reg_ram_208__6 (.Q (camera_module_cache_ram_208__6)
         , .QB (\$dummy [40]), .D (nx19103), .CLK (clk), .R (rst)) ;
    mux21_ni ix19104 (.Y (nx19103), .A0 (camera_module_cache_ram_208__6), .A1 (
             nx35522), .S0 (nx35082)) ;
    aoi22 ix23283 (.Y (nx23282), .A0 (camera_module_cache_ram_224__6), .A1 (
          nx36368), .B0 (camera_module_cache_ram_240__6), .B1 (nx36408)) ;
    dffr camera_module_cache_reg_ram_224__6 (.Q (camera_module_cache_ram_224__6)
         , .QB (\$dummy [41]), .D (nx19093), .CLK (clk), .R (rst)) ;
    mux21_ni ix19094 (.Y (nx19093), .A0 (camera_module_cache_ram_224__6), .A1 (
             nx35524), .S0 (nx35078)) ;
    dffr camera_module_cache_reg_ram_240__6 (.Q (camera_module_cache_ram_240__6)
         , .QB (\$dummy [42]), .D (nx19083), .CLK (clk), .R (rst)) ;
    mux21_ni ix19084 (.Y (nx19083), .A0 (camera_module_cache_ram_240__6), .A1 (
             nx35524), .S0 (nx35074)) ;
    nor02_2x ix23299 (.Y (nx23298), .A0 (nx1056), .A1 (nx986)) ;
    oai21 ix23303 (.Y (nx23302), .A0 (nx22416), .A1 (nx22338), .B0 (nx36452)) ;
    nand04 ix22417 (.Y (nx22416), .A0 (nx23305), .A1 (nx23324), .A2 (nx23337), .A3 (
           nx23349)) ;
    aoi22 ix23306 (.Y (nx23305), .A0 (camera_module_cache_ram_1__6), .A1 (
          nx37030), .B0 (camera_module_cache_ram_17__6), .B1 (nx37032)) ;
    dffr camera_module_cache_reg_ram_1__6 (.Q (camera_module_cache_ram_1__6), .QB (
         \$dummy [43]), .D (nx19073), .CLK (clk), .R (rst)) ;
    mux21_ni ix19074 (.Y (nx19073), .A0 (camera_module_cache_ram_1__6), .A1 (
             nx35524), .S0 (nx35064)) ;
    nand02 ix5359 (.Y (nx5358), .A0 (nx23314), .A1 (nx23091)) ;
    dffr camera_module_cache_reg_ram_17__6 (.Q (camera_module_cache_ram_17__6), 
         .QB (\$dummy [44]), .D (nx19063), .CLK (clk), .R (rst)) ;
    mux21_ni ix19064 (.Y (nx19063), .A0 (camera_module_cache_ram_17__6), .A1 (
             nx35524), .S0 (nx35060)) ;
    aoi22 ix23325 (.Y (nx23324), .A0 (camera_module_cache_ram_33__6), .A1 (
          nx37034), .B0 (camera_module_cache_ram_49__6), .B1 (nx37036)) ;
    dffr camera_module_cache_reg_ram_33__6 (.Q (camera_module_cache_ram_33__6), 
         .QB (\$dummy [45]), .D (nx19053), .CLK (clk), .R (rst)) ;
    mux21_ni ix19054 (.Y (nx19053), .A0 (camera_module_cache_ram_33__6), .A1 (
             nx35524), .S0 (nx35056)) ;
    dffr camera_module_cache_reg_ram_49__6 (.Q (camera_module_cache_ram_49__6), 
         .QB (\$dummy [46]), .D (nx19043), .CLK (clk), .R (rst)) ;
    mux21_ni ix19044 (.Y (nx19043), .A0 (camera_module_cache_ram_49__6), .A1 (
             nx35524), .S0 (nx35052)) ;
    aoi22 ix23338 (.Y (nx23337), .A0 (camera_module_cache_ram_65__6), .A1 (
          nx37038), .B0 (camera_module_cache_ram_81__6), .B1 (nx37040)) ;
    dffr camera_module_cache_reg_ram_65__6 (.Q (camera_module_cache_ram_65__6), 
         .QB (\$dummy [47]), .D (nx19033), .CLK (clk), .R (rst)) ;
    mux21_ni ix19034 (.Y (nx19033), .A0 (camera_module_cache_ram_65__6), .A1 (
             nx35524), .S0 (nx35048)) ;
    dffr camera_module_cache_reg_ram_81__6 (.Q (camera_module_cache_ram_81__6), 
         .QB (\$dummy [48]), .D (nx19023), .CLK (clk), .R (rst)) ;
    mux21_ni ix19024 (.Y (nx19023), .A0 (camera_module_cache_ram_81__6), .A1 (
             nx35526), .S0 (nx35044)) ;
    aoi22 ix23350 (.Y (nx23349), .A0 (camera_module_cache_ram_113__6), .A1 (
          nx37042), .B0 (camera_module_cache_ram_97__6), .B1 (nx37044)) ;
    dffr camera_module_cache_reg_ram_113__6 (.Q (camera_module_cache_ram_113__6)
         , .QB (\$dummy [49]), .D (nx19003), .CLK (clk), .R (rst)) ;
    mux21_ni ix19004 (.Y (nx19003), .A0 (camera_module_cache_ram_113__6), .A1 (
             nx35526), .S0 (nx35036)) ;
    dffr camera_module_cache_reg_ram_97__6 (.Q (camera_module_cache_ram_97__6), 
         .QB (\$dummy [50]), .D (nx19013), .CLK (clk), .R (rst)) ;
    mux21_ni ix19014 (.Y (nx19013), .A0 (camera_module_cache_ram_97__6), .A1 (
             nx35526), .S0 (nx35040)) ;
    nand04 ix22339 (.Y (nx22338), .A0 (nx23361), .A1 (nx23372), .A2 (nx23385), .A3 (
           nx23400)) ;
    aoi22 ix23362 (.Y (nx23361), .A0 (camera_module_cache_ram_129__6), .A1 (
          nx37046), .B0 (camera_module_cache_ram_145__6), .B1 (nx37048)) ;
    dffr camera_module_cache_reg_ram_129__6 (.Q (camera_module_cache_ram_129__6)
         , .QB (\$dummy [51]), .D (nx18993), .CLK (clk), .R (rst)) ;
    mux21_ni ix18994 (.Y (nx18993), .A0 (camera_module_cache_ram_129__6), .A1 (
             nx35526), .S0 (nx35032)) ;
    dffr camera_module_cache_reg_ram_145__6 (.Q (camera_module_cache_ram_145__6)
         , .QB (\$dummy [52]), .D (nx18983), .CLK (clk), .R (rst)) ;
    mux21_ni ix18984 (.Y (nx18983), .A0 (camera_module_cache_ram_145__6), .A1 (
             nx35526), .S0 (nx35028)) ;
    aoi22 ix23373 (.Y (nx23372), .A0 (camera_module_cache_ram_177__6), .A1 (
          nx37050), .B0 (camera_module_cache_ram_161__6), .B1 (nx37052)) ;
    dffr camera_module_cache_reg_ram_177__6 (.Q (camera_module_cache_ram_177__6)
         , .QB (\$dummy [53]), .D (nx18963), .CLK (clk), .R (rst)) ;
    mux21_ni ix18964 (.Y (nx18963), .A0 (camera_module_cache_ram_177__6), .A1 (
             nx35526), .S0 (nx35020)) ;
    dffr camera_module_cache_reg_ram_161__6 (.Q (camera_module_cache_ram_161__6)
         , .QB (\$dummy [54]), .D (nx18973), .CLK (clk), .R (rst)) ;
    mux21_ni ix18974 (.Y (nx18973), .A0 (camera_module_cache_ram_161__6), .A1 (
             nx35526), .S0 (nx35024)) ;
    aoi22 ix23386 (.Y (nx23385), .A0 (camera_module_cache_ram_193__6), .A1 (
          nx36288), .B0 (camera_module_cache_ram_209__6), .B1 (nx36328)) ;
    dffr camera_module_cache_reg_ram_193__6 (.Q (camera_module_cache_ram_193__6)
         , .QB (\$dummy [55]), .D (nx18953), .CLK (clk), .R (rst)) ;
    mux21_ni ix18954 (.Y (nx18953), .A0 (camera_module_cache_ram_193__6), .A1 (
             nx35528), .S0 (nx35016)) ;
    dffr camera_module_cache_reg_ram_209__6 (.Q (camera_module_cache_ram_209__6)
         , .QB (\$dummy [56]), .D (nx18943), .CLK (clk), .R (rst)) ;
    mux21_ni ix18944 (.Y (nx18943), .A0 (camera_module_cache_ram_209__6), .A1 (
             nx35528), .S0 (nx35012)) ;
    aoi22 ix23401 (.Y (nx23400), .A0 (camera_module_cache_ram_225__6), .A1 (
          nx36368), .B0 (camera_module_cache_ram_241__6), .B1 (nx36408)) ;
    dffr camera_module_cache_reg_ram_225__6 (.Q (camera_module_cache_ram_225__6)
         , .QB (\$dummy [57]), .D (nx18933), .CLK (clk), .R (rst)) ;
    mux21_ni ix18934 (.Y (nx18933), .A0 (camera_module_cache_ram_225__6), .A1 (
             nx35528), .S0 (nx35008)) ;
    dffr camera_module_cache_reg_ram_241__6 (.Q (camera_module_cache_ram_241__6)
         , .QB (\$dummy [58]), .D (nx18923), .CLK (clk), .R (rst)) ;
    mux21_ni ix18924 (.Y (nx18923), .A0 (camera_module_cache_ram_241__6), .A1 (
             nx35528), .S0 (nx35004)) ;
    oai21 ix23414 (.Y (nx23413), .A0 (nx22252), .A1 (nx22174), .B0 (nx36456)) ;
    nand04 ix22253 (.Y (nx22252), .A0 (nx23417), .A1 (nx23433), .A2 (nx23446), .A3 (
           nx23458)) ;
    aoi22 ix23418 (.Y (nx23417), .A0 (camera_module_cache_ram_2__6), .A1 (
          nx37030), .B0 (camera_module_cache_ram_18__6), .B1 (nx37032)) ;
    dffr camera_module_cache_reg_ram_2__6 (.Q (camera_module_cache_ram_2__6), .QB (
         \$dummy [59]), .D (nx18913), .CLK (clk), .R (rst)) ;
    mux21_ni ix18914 (.Y (nx18913), .A0 (camera_module_cache_ram_2__6), .A1 (
             nx35528), .S0 (nx34994)) ;
    nand02 ix5065 (.Y (nx5064), .A0 (nx23423), .A1 (nx23091)) ;
    dffr camera_module_cache_reg_ram_18__6 (.Q (camera_module_cache_ram_18__6), 
         .QB (\$dummy [60]), .D (nx18903), .CLK (clk), .R (rst)) ;
    mux21_ni ix18904 (.Y (nx18903), .A0 (camera_module_cache_ram_18__6), .A1 (
             nx35528), .S0 (nx34990)) ;
    aoi22 ix23434 (.Y (nx23433), .A0 (camera_module_cache_ram_34__6), .A1 (
          nx37034), .B0 (camera_module_cache_ram_50__6), .B1 (nx37036)) ;
    dffr camera_module_cache_reg_ram_34__6 (.Q (camera_module_cache_ram_34__6), 
         .QB (\$dummy [61]), .D (nx18893), .CLK (clk), .R (rst)) ;
    mux21_ni ix18894 (.Y (nx18893), .A0 (camera_module_cache_ram_34__6), .A1 (
             nx35528), .S0 (nx34986)) ;
    dffr camera_module_cache_reg_ram_50__6 (.Q (camera_module_cache_ram_50__6), 
         .QB (\$dummy [62]), .D (nx18883), .CLK (clk), .R (rst)) ;
    mux21_ni ix18884 (.Y (nx18883), .A0 (camera_module_cache_ram_50__6), .A1 (
             nx35530), .S0 (nx34982)) ;
    aoi22 ix23447 (.Y (nx23446), .A0 (camera_module_cache_ram_66__6), .A1 (
          nx37038), .B0 (camera_module_cache_ram_82__6), .B1 (nx37040)) ;
    dffr camera_module_cache_reg_ram_66__6 (.Q (camera_module_cache_ram_66__6), 
         .QB (\$dummy [63]), .D (nx18873), .CLK (clk), .R (rst)) ;
    mux21_ni ix18874 (.Y (nx18873), .A0 (camera_module_cache_ram_66__6), .A1 (
             nx35530), .S0 (nx34978)) ;
    dffr camera_module_cache_reg_ram_82__6 (.Q (camera_module_cache_ram_82__6), 
         .QB (\$dummy [64]), .D (nx18863), .CLK (clk), .R (rst)) ;
    mux21_ni ix18864 (.Y (nx18863), .A0 (camera_module_cache_ram_82__6), .A1 (
             nx35530), .S0 (nx34974)) ;
    aoi22 ix23459 (.Y (nx23458), .A0 (camera_module_cache_ram_114__6), .A1 (
          nx37042), .B0 (camera_module_cache_ram_98__6), .B1 (nx37044)) ;
    dffr camera_module_cache_reg_ram_114__6 (.Q (camera_module_cache_ram_114__6)
         , .QB (\$dummy [65]), .D (nx18843), .CLK (clk), .R (rst)) ;
    mux21_ni ix18844 (.Y (nx18843), .A0 (camera_module_cache_ram_114__6), .A1 (
             nx35530), .S0 (nx34966)) ;
    dffr camera_module_cache_reg_ram_98__6 (.Q (camera_module_cache_ram_98__6), 
         .QB (\$dummy [66]), .D (nx18853), .CLK (clk), .R (rst)) ;
    mux21_ni ix18854 (.Y (nx18853), .A0 (camera_module_cache_ram_98__6), .A1 (
             nx35530), .S0 (nx34970)) ;
    nand04 ix22175 (.Y (nx22174), .A0 (nx23469), .A1 (nx23482), .A2 (nx23495), .A3 (
           nx23506)) ;
    aoi22 ix23470 (.Y (nx23469), .A0 (camera_module_cache_ram_130__6), .A1 (
          nx37046), .B0 (camera_module_cache_ram_146__6), .B1 (nx37048)) ;
    dffr camera_module_cache_reg_ram_130__6 (.Q (camera_module_cache_ram_130__6)
         , .QB (\$dummy [67]), .D (nx18833), .CLK (clk), .R (rst)) ;
    mux21_ni ix18834 (.Y (nx18833), .A0 (camera_module_cache_ram_130__6), .A1 (
             nx35530), .S0 (nx34962)) ;
    dffr camera_module_cache_reg_ram_146__6 (.Q (camera_module_cache_ram_146__6)
         , .QB (\$dummy [68]), .D (nx18823), .CLK (clk), .R (rst)) ;
    mux21_ni ix18824 (.Y (nx18823), .A0 (camera_module_cache_ram_146__6), .A1 (
             nx35530), .S0 (nx34958)) ;
    aoi22 ix23483 (.Y (nx23482), .A0 (camera_module_cache_ram_178__6), .A1 (
          nx37050), .B0 (camera_module_cache_ram_162__6), .B1 (nx37052)) ;
    dffr camera_module_cache_reg_ram_178__6 (.Q (camera_module_cache_ram_178__6)
         , .QB (\$dummy [69]), .D (nx18803), .CLK (clk), .R (rst)) ;
    mux21_ni ix18804 (.Y (nx18803), .A0 (camera_module_cache_ram_178__6), .A1 (
             nx35532), .S0 (nx34950)) ;
    dffr camera_module_cache_reg_ram_162__6 (.Q (camera_module_cache_ram_162__6)
         , .QB (\$dummy [70]), .D (nx18813), .CLK (clk), .R (rst)) ;
    mux21_ni ix18814 (.Y (nx18813), .A0 (camera_module_cache_ram_162__6), .A1 (
             nx35532), .S0 (nx34954)) ;
    aoi22 ix23496 (.Y (nx23495), .A0 (camera_module_cache_ram_194__6), .A1 (
          nx36288), .B0 (camera_module_cache_ram_210__6), .B1 (nx36328)) ;
    dffr camera_module_cache_reg_ram_194__6 (.Q (camera_module_cache_ram_194__6)
         , .QB (\$dummy [71]), .D (nx18793), .CLK (clk), .R (rst)) ;
    mux21_ni ix18794 (.Y (nx18793), .A0 (camera_module_cache_ram_194__6), .A1 (
             nx35532), .S0 (nx34946)) ;
    dffr camera_module_cache_reg_ram_210__6 (.Q (camera_module_cache_ram_210__6)
         , .QB (\$dummy [72]), .D (nx18783), .CLK (clk), .R (rst)) ;
    mux21_ni ix18784 (.Y (nx18783), .A0 (camera_module_cache_ram_210__6), .A1 (
             nx35532), .S0 (nx34942)) ;
    aoi22 ix23507 (.Y (nx23506), .A0 (camera_module_cache_ram_226__6), .A1 (
          nx36368), .B0 (camera_module_cache_ram_242__6), .B1 (nx36408)) ;
    dffr camera_module_cache_reg_ram_226__6 (.Q (camera_module_cache_ram_226__6)
         , .QB (\$dummy [73]), .D (nx18773), .CLK (clk), .R (rst)) ;
    mux21_ni ix18774 (.Y (nx18773), .A0 (camera_module_cache_ram_226__6), .A1 (
             nx35532), .S0 (nx34938)) ;
    dffr camera_module_cache_reg_ram_242__6 (.Q (camera_module_cache_ram_242__6)
         , .QB (\$dummy [74]), .D (nx18763), .CLK (clk), .R (rst)) ;
    mux21_ni ix18764 (.Y (nx18763), .A0 (camera_module_cache_ram_242__6), .A1 (
             nx35532), .S0 (nx34934)) ;
    oai21 ix23521 (.Y (nx23520), .A0 (nx22090), .A1 (nx22012), .B0 (nx36460)) ;
    nand04 ix22091 (.Y (nx22090), .A0 (nx23523), .A1 (nx23537), .A2 (nx23549), .A3 (
           nx23562)) ;
    aoi22 ix23524 (.Y (nx23523), .A0 (camera_module_cache_ram_3__6), .A1 (
          nx37030), .B0 (camera_module_cache_ram_19__6), .B1 (nx37032)) ;
    dffr camera_module_cache_reg_ram_3__6 (.Q (camera_module_cache_ram_3__6), .QB (
         \$dummy [75]), .D (nx18753), .CLK (clk), .R (rst)) ;
    mux21_ni ix18754 (.Y (nx18753), .A0 (camera_module_cache_ram_3__6), .A1 (
             nx35532), .S0 (nx34924)) ;
    nand02 ix4773 (.Y (nx4772), .A0 (nx23529), .A1 (nx23091)) ;
    dffr camera_module_cache_reg_ram_19__6 (.Q (camera_module_cache_ram_19__6), 
         .QB (\$dummy [76]), .D (nx18743), .CLK (clk), .R (rst)) ;
    mux21_ni ix18744 (.Y (nx18743), .A0 (camera_module_cache_ram_19__6), .A1 (
             nx35534), .S0 (nx34920)) ;
    aoi22 ix23538 (.Y (nx23537), .A0 (camera_module_cache_ram_35__6), .A1 (
          nx37034), .B0 (camera_module_cache_ram_51__6), .B1 (nx37036)) ;
    dffr camera_module_cache_reg_ram_35__6 (.Q (camera_module_cache_ram_35__6), 
         .QB (\$dummy [77]), .D (nx18733), .CLK (clk), .R (rst)) ;
    mux21_ni ix18734 (.Y (nx18733), .A0 (camera_module_cache_ram_35__6), .A1 (
             nx35534), .S0 (nx34916)) ;
    dffr camera_module_cache_reg_ram_51__6 (.Q (camera_module_cache_ram_51__6), 
         .QB (\$dummy [78]), .D (nx18723), .CLK (clk), .R (rst)) ;
    mux21_ni ix18724 (.Y (nx18723), .A0 (camera_module_cache_ram_51__6), .A1 (
             nx35534), .S0 (nx34912)) ;
    aoi22 ix23550 (.Y (nx23549), .A0 (camera_module_cache_ram_67__6), .A1 (
          nx37038), .B0 (camera_module_cache_ram_83__6), .B1 (nx37040)) ;
    dffr camera_module_cache_reg_ram_67__6 (.Q (camera_module_cache_ram_67__6), 
         .QB (\$dummy [79]), .D (nx18713), .CLK (clk), .R (rst)) ;
    mux21_ni ix18714 (.Y (nx18713), .A0 (camera_module_cache_ram_67__6), .A1 (
             nx35534), .S0 (nx34908)) ;
    dffr camera_module_cache_reg_ram_83__6 (.Q (camera_module_cache_ram_83__6), 
         .QB (\$dummy [80]), .D (nx18703), .CLK (clk), .R (rst)) ;
    mux21_ni ix18704 (.Y (nx18703), .A0 (camera_module_cache_ram_83__6), .A1 (
             nx35534), .S0 (nx34904)) ;
    aoi22 ix23563 (.Y (nx23562), .A0 (camera_module_cache_ram_115__6), .A1 (
          nx37042), .B0 (camera_module_cache_ram_99__6), .B1 (nx37044)) ;
    dffr camera_module_cache_reg_ram_115__6 (.Q (camera_module_cache_ram_115__6)
         , .QB (\$dummy [81]), .D (nx18683), .CLK (clk), .R (rst)) ;
    mux21_ni ix18684 (.Y (nx18683), .A0 (camera_module_cache_ram_115__6), .A1 (
             nx35534), .S0 (nx34896)) ;
    dffr camera_module_cache_reg_ram_99__6 (.Q (camera_module_cache_ram_99__6), 
         .QB (\$dummy [82]), .D (nx18693), .CLK (clk), .R (rst)) ;
    mux21_ni ix18694 (.Y (nx18693), .A0 (camera_module_cache_ram_99__6), .A1 (
             nx35534), .S0 (nx34900)) ;
    nand04 ix22013 (.Y (nx22012), .A0 (nx23574), .A1 (nx23587), .A2 (nx23599), .A3 (
           nx23610)) ;
    aoi22 ix23575 (.Y (nx23574), .A0 (camera_module_cache_ram_131__6), .A1 (
          nx37046), .B0 (camera_module_cache_ram_147__6), .B1 (nx37048)) ;
    dffr camera_module_cache_reg_ram_131__6 (.Q (camera_module_cache_ram_131__6)
         , .QB (\$dummy [83]), .D (nx18673), .CLK (clk), .R (rst)) ;
    mux21_ni ix18674 (.Y (nx18673), .A0 (camera_module_cache_ram_131__6), .A1 (
             nx35536), .S0 (nx34892)) ;
    dffr camera_module_cache_reg_ram_147__6 (.Q (camera_module_cache_ram_147__6)
         , .QB (\$dummy [84]), .D (nx18663), .CLK (clk), .R (rst)) ;
    mux21_ni ix18664 (.Y (nx18663), .A0 (camera_module_cache_ram_147__6), .A1 (
             nx35536), .S0 (nx34888)) ;
    aoi22 ix23588 (.Y (nx23587), .A0 (camera_module_cache_ram_179__6), .A1 (
          nx37050), .B0 (camera_module_cache_ram_163__6), .B1 (nx37052)) ;
    dffr camera_module_cache_reg_ram_179__6 (.Q (camera_module_cache_ram_179__6)
         , .QB (\$dummy [85]), .D (nx18643), .CLK (clk), .R (rst)) ;
    mux21_ni ix18644 (.Y (nx18643), .A0 (camera_module_cache_ram_179__6), .A1 (
             nx35536), .S0 (nx34880)) ;
    dffr camera_module_cache_reg_ram_163__6 (.Q (camera_module_cache_ram_163__6)
         , .QB (\$dummy [86]), .D (nx18653), .CLK (clk), .R (rst)) ;
    mux21_ni ix18654 (.Y (nx18653), .A0 (camera_module_cache_ram_163__6), .A1 (
             nx35536), .S0 (nx34884)) ;
    aoi22 ix23600 (.Y (nx23599), .A0 (camera_module_cache_ram_195__6), .A1 (
          nx36288), .B0 (camera_module_cache_ram_211__6), .B1 (nx36328)) ;
    dffr camera_module_cache_reg_ram_195__6 (.Q (camera_module_cache_ram_195__6)
         , .QB (\$dummy [87]), .D (nx18633), .CLK (clk), .R (rst)) ;
    mux21_ni ix18634 (.Y (nx18633), .A0 (camera_module_cache_ram_195__6), .A1 (
             nx35536), .S0 (nx34876)) ;
    dffr camera_module_cache_reg_ram_211__6 (.Q (camera_module_cache_ram_211__6)
         , .QB (\$dummy [88]), .D (nx18623), .CLK (clk), .R (rst)) ;
    mux21_ni ix18624 (.Y (nx18623), .A0 (camera_module_cache_ram_211__6), .A1 (
             nx35536), .S0 (nx34872)) ;
    aoi22 ix23611 (.Y (nx23610), .A0 (camera_module_cache_ram_227__6), .A1 (
          nx36368), .B0 (camera_module_cache_ram_243__6), .B1 (nx36408)) ;
    dffr camera_module_cache_reg_ram_227__6 (.Q (camera_module_cache_ram_227__6)
         , .QB (\$dummy [89]), .D (nx18613), .CLK (clk), .R (rst)) ;
    mux21_ni ix18614 (.Y (nx18613), .A0 (camera_module_cache_ram_227__6), .A1 (
             nx35536), .S0 (nx34868)) ;
    dffr camera_module_cache_reg_ram_243__6 (.Q (camera_module_cache_ram_243__6)
         , .QB (\$dummy [90]), .D (nx18603), .CLK (clk), .R (rst)) ;
    mux21_ni ix18604 (.Y (nx18603), .A0 (camera_module_cache_ram_243__6), .A1 (
             nx35538), .S0 (nx34864)) ;
    nand02 ix843 (.Y (nx842), .A0 (nx836), .A1 (nx810)) ;
    nand04 ix21935 (.Y (nx21934), .A0 (nx23627), .A1 (nx23733), .A2 (nx23835), .A3 (
           nx23938)) ;
    oai21 ix23628 (.Y (nx23627), .A0 (nx21924), .A1 (nx21846), .B0 (nx36464)) ;
    nand04 ix21925 (.Y (nx21924), .A0 (nx23630), .A1 (nx23648), .A2 (nx23660), .A3 (
           nx23670)) ;
    aoi22 ix23631 (.Y (nx23630), .A0 (camera_module_cache_ram_4__6), .A1 (
          nx37030), .B0 (camera_module_cache_ram_20__6), .B1 (nx37032)) ;
    dffr camera_module_cache_reg_ram_4__6 (.Q (camera_module_cache_ram_4__6), .QB (
         \$dummy [91]), .D (nx18593), .CLK (clk), .R (rst)) ;
    mux21_ni ix18594 (.Y (nx18593), .A0 (camera_module_cache_ram_4__6), .A1 (
             nx35538), .S0 (nx34854)) ;
    nand02 ix4475 (.Y (nx4474), .A0 (nx23639), .A1 (nx23105)) ;
    dffr camera_module_cache_reg_ram_20__6 (.Q (camera_module_cache_ram_20__6), 
         .QB (\$dummy [92]), .D (nx18583), .CLK (clk), .R (rst)) ;
    mux21_ni ix18584 (.Y (nx18583), .A0 (camera_module_cache_ram_20__6), .A1 (
             nx35538), .S0 (nx34850)) ;
    aoi22 ix23649 (.Y (nx23648), .A0 (camera_module_cache_ram_36__6), .A1 (
          nx37034), .B0 (camera_module_cache_ram_52__6), .B1 (nx37036)) ;
    dffr camera_module_cache_reg_ram_36__6 (.Q (camera_module_cache_ram_36__6), 
         .QB (\$dummy [93]), .D (nx18573), .CLK (clk), .R (rst)) ;
    mux21_ni ix18574 (.Y (nx18573), .A0 (camera_module_cache_ram_36__6), .A1 (
             nx35538), .S0 (nx34846)) ;
    dffr camera_module_cache_reg_ram_52__6 (.Q (camera_module_cache_ram_52__6), 
         .QB (\$dummy [94]), .D (nx18563), .CLK (clk), .R (rst)) ;
    mux21_ni ix18564 (.Y (nx18563), .A0 (camera_module_cache_ram_52__6), .A1 (
             nx35538), .S0 (nx34842)) ;
    aoi22 ix23661 (.Y (nx23660), .A0 (camera_module_cache_ram_68__6), .A1 (
          nx37038), .B0 (camera_module_cache_ram_84__6), .B1 (nx37040)) ;
    dffr camera_module_cache_reg_ram_68__6 (.Q (camera_module_cache_ram_68__6), 
         .QB (\$dummy [95]), .D (nx18553), .CLK (clk), .R (rst)) ;
    mux21_ni ix18554 (.Y (nx18553), .A0 (camera_module_cache_ram_68__6), .A1 (
             nx35538), .S0 (nx34838)) ;
    dffr camera_module_cache_reg_ram_84__6 (.Q (camera_module_cache_ram_84__6), 
         .QB (\$dummy [96]), .D (nx18543), .CLK (clk), .R (rst)) ;
    mux21_ni ix18544 (.Y (nx18543), .A0 (camera_module_cache_ram_84__6), .A1 (
             nx35538), .S0 (nx34834)) ;
    aoi22 ix23671 (.Y (nx23670), .A0 (camera_module_cache_ram_116__6), .A1 (
          nx37042), .B0 (camera_module_cache_ram_100__6), .B1 (nx37044)) ;
    dffr camera_module_cache_reg_ram_116__6 (.Q (camera_module_cache_ram_116__6)
         , .QB (\$dummy [97]), .D (nx18523), .CLK (clk), .R (rst)) ;
    mux21_ni ix18524 (.Y (nx18523), .A0 (camera_module_cache_ram_116__6), .A1 (
             nx35540), .S0 (nx34826)) ;
    dffr camera_module_cache_reg_ram_100__6 (.Q (camera_module_cache_ram_100__6)
         , .QB (\$dummy [98]), .D (nx18533), .CLK (clk), .R (rst)) ;
    mux21_ni ix18534 (.Y (nx18533), .A0 (camera_module_cache_ram_100__6), .A1 (
             nx35540), .S0 (nx34830)) ;
    nand04 ix21847 (.Y (nx21846), .A0 (nx23683), .A1 (nx23695), .A2 (nx23706), .A3 (
           nx23719)) ;
    aoi22 ix23684 (.Y (nx23683), .A0 (camera_module_cache_ram_132__6), .A1 (
          nx37046), .B0 (camera_module_cache_ram_148__6), .B1 (nx37048)) ;
    dffr camera_module_cache_reg_ram_132__6 (.Q (camera_module_cache_ram_132__6)
         , .QB (\$dummy [99]), .D (nx18513), .CLK (clk), .R (rst)) ;
    mux21_ni ix18514 (.Y (nx18513), .A0 (camera_module_cache_ram_132__6), .A1 (
             nx35540), .S0 (nx34822)) ;
    dffr camera_module_cache_reg_ram_148__6 (.Q (camera_module_cache_ram_148__6)
         , .QB (\$dummy [100]), .D (nx18503), .CLK (clk), .R (rst)) ;
    mux21_ni ix18504 (.Y (nx18503), .A0 (camera_module_cache_ram_148__6), .A1 (
             nx35540), .S0 (nx34818)) ;
    aoi22 ix23696 (.Y (nx23695), .A0 (camera_module_cache_ram_180__6), .A1 (
          nx37050), .B0 (camera_module_cache_ram_164__6), .B1 (nx37052)) ;
    dffr camera_module_cache_reg_ram_180__6 (.Q (camera_module_cache_ram_180__6)
         , .QB (\$dummy [101]), .D (nx18483), .CLK (clk), .R (rst)) ;
    mux21_ni ix18484 (.Y (nx18483), .A0 (camera_module_cache_ram_180__6), .A1 (
             nx35540), .S0 (nx34810)) ;
    dffr camera_module_cache_reg_ram_164__6 (.Q (camera_module_cache_ram_164__6)
         , .QB (\$dummy [102]), .D (nx18493), .CLK (clk), .R (rst)) ;
    mux21_ni ix18494 (.Y (nx18493), .A0 (camera_module_cache_ram_164__6), .A1 (
             nx35540), .S0 (nx34814)) ;
    aoi22 ix23707 (.Y (nx23706), .A0 (camera_module_cache_ram_196__6), .A1 (
          nx36288), .B0 (camera_module_cache_ram_212__6), .B1 (nx36328)) ;
    dffr camera_module_cache_reg_ram_196__6 (.Q (camera_module_cache_ram_196__6)
         , .QB (\$dummy [103]), .D (nx18473), .CLK (clk), .R (rst)) ;
    mux21_ni ix18474 (.Y (nx18473), .A0 (camera_module_cache_ram_196__6), .A1 (
             nx35540), .S0 (nx34806)) ;
    dffr camera_module_cache_reg_ram_212__6 (.Q (camera_module_cache_ram_212__6)
         , .QB (\$dummy [104]), .D (nx18463), .CLK (clk), .R (rst)) ;
    mux21_ni ix18464 (.Y (nx18463), .A0 (camera_module_cache_ram_212__6), .A1 (
             nx35542), .S0 (nx34802)) ;
    aoi22 ix23720 (.Y (nx23719), .A0 (camera_module_cache_ram_228__6), .A1 (
          nx36368), .B0 (camera_module_cache_ram_244__6), .B1 (nx36408)) ;
    dffr camera_module_cache_reg_ram_228__6 (.Q (camera_module_cache_ram_228__6)
         , .QB (\$dummy [105]), .D (nx18453), .CLK (clk), .R (rst)) ;
    mux21_ni ix18454 (.Y (nx18453), .A0 (camera_module_cache_ram_228__6), .A1 (
             nx35542), .S0 (nx34798)) ;
    dffr camera_module_cache_reg_ram_244__6 (.Q (camera_module_cache_ram_244__6)
         , .QB (\$dummy [106]), .D (nx18443), .CLK (clk), .R (rst)) ;
    mux21_ni ix18444 (.Y (nx18443), .A0 (camera_module_cache_ram_244__6), .A1 (
             nx35542), .S0 (nx34794)) ;
    oai21 ix23734 (.Y (nx23733), .A0 (nx21762), .A1 (nx21684), .B0 (nx36468)) ;
    nand04 ix21763 (.Y (nx21762), .A0 (nx23736), .A1 (nx23748), .A2 (nx23761), .A3 (
           nx23772)) ;
    aoi22 ix23737 (.Y (nx23736), .A0 (camera_module_cache_ram_5__6), .A1 (
          nx37030), .B0 (camera_module_cache_ram_21__6), .B1 (nx37032)) ;
    dffr camera_module_cache_reg_ram_5__6 (.Q (camera_module_cache_ram_5__6), .QB (
         \$dummy [107]), .D (nx18433), .CLK (clk), .R (rst)) ;
    mux21_ni ix18434 (.Y (nx18433), .A0 (camera_module_cache_ram_5__6), .A1 (
             nx35542), .S0 (nx34784)) ;
    nand02 ix4183 (.Y (nx4182), .A0 (nx23639), .A1 (nx23314)) ;
    dffr camera_module_cache_reg_ram_21__6 (.Q (camera_module_cache_ram_21__6), 
         .QB (\$dummy [108]), .D (nx18423), .CLK (clk), .R (rst)) ;
    mux21_ni ix18424 (.Y (nx18423), .A0 (camera_module_cache_ram_21__6), .A1 (
             nx35542), .S0 (nx34780)) ;
    aoi22 ix23749 (.Y (nx23748), .A0 (camera_module_cache_ram_37__6), .A1 (
          nx37034), .B0 (camera_module_cache_ram_53__6), .B1 (nx37036)) ;
    dffr camera_module_cache_reg_ram_37__6 (.Q (camera_module_cache_ram_37__6), 
         .QB (\$dummy [109]), .D (nx18413), .CLK (clk), .R (rst)) ;
    mux21_ni ix18414 (.Y (nx18413), .A0 (camera_module_cache_ram_37__6), .A1 (
             nx35542), .S0 (nx34776)) ;
    dffr camera_module_cache_reg_ram_53__6 (.Q (camera_module_cache_ram_53__6), 
         .QB (\$dummy [110]), .D (nx18403), .CLK (clk), .R (rst)) ;
    mux21_ni ix18404 (.Y (nx18403), .A0 (camera_module_cache_ram_53__6), .A1 (
             nx35542), .S0 (nx34772)) ;
    aoi22 ix23762 (.Y (nx23761), .A0 (camera_module_cache_ram_69__6), .A1 (
          nx37038), .B0 (camera_module_cache_ram_85__6), .B1 (nx37040)) ;
    dffr camera_module_cache_reg_ram_69__6 (.Q (camera_module_cache_ram_69__6), 
         .QB (\$dummy [111]), .D (nx18393), .CLK (clk), .R (rst)) ;
    mux21_ni ix18394 (.Y (nx18393), .A0 (camera_module_cache_ram_69__6), .A1 (
             nx35544), .S0 (nx34768)) ;
    dffr camera_module_cache_reg_ram_85__6 (.Q (camera_module_cache_ram_85__6), 
         .QB (\$dummy [112]), .D (nx18383), .CLK (clk), .R (rst)) ;
    mux21_ni ix18384 (.Y (nx18383), .A0 (camera_module_cache_ram_85__6), .A1 (
             nx35544), .S0 (nx34764)) ;
    aoi22 ix23773 (.Y (nx23772), .A0 (camera_module_cache_ram_117__6), .A1 (
          nx37042), .B0 (camera_module_cache_ram_101__6), .B1 (nx37044)) ;
    dffr camera_module_cache_reg_ram_117__6 (.Q (camera_module_cache_ram_117__6)
         , .QB (\$dummy [113]), .D (nx18363), .CLK (clk), .R (rst)) ;
    mux21_ni ix18364 (.Y (nx18363), .A0 (camera_module_cache_ram_117__6), .A1 (
             nx35544), .S0 (nx34756)) ;
    dffr camera_module_cache_reg_ram_101__6 (.Q (camera_module_cache_ram_101__6)
         , .QB (\$dummy [114]), .D (nx18373), .CLK (clk), .R (rst)) ;
    mux21_ni ix18374 (.Y (nx18373), .A0 (camera_module_cache_ram_101__6), .A1 (
             nx35544), .S0 (nx34760)) ;
    nand04 ix21685 (.Y (nx21684), .A0 (nx23785), .A1 (nx23797), .A2 (nx23811), .A3 (
           nx23822)) ;
    aoi22 ix23786 (.Y (nx23785), .A0 (camera_module_cache_ram_133__6), .A1 (
          nx37046), .B0 (camera_module_cache_ram_149__6), .B1 (nx37048)) ;
    dffr camera_module_cache_reg_ram_133__6 (.Q (camera_module_cache_ram_133__6)
         , .QB (\$dummy [115]), .D (nx18353), .CLK (clk), .R (rst)) ;
    mux21_ni ix18354 (.Y (nx18353), .A0 (camera_module_cache_ram_133__6), .A1 (
             nx35544), .S0 (nx34752)) ;
    dffr camera_module_cache_reg_ram_149__6 (.Q (camera_module_cache_ram_149__6)
         , .QB (\$dummy [116]), .D (nx18343), .CLK (clk), .R (rst)) ;
    mux21_ni ix18344 (.Y (nx18343), .A0 (camera_module_cache_ram_149__6), .A1 (
             nx35544), .S0 (nx34748)) ;
    aoi22 ix23798 (.Y (nx23797), .A0 (camera_module_cache_ram_181__6), .A1 (
          nx37050), .B0 (camera_module_cache_ram_165__6), .B1 (nx37052)) ;
    dffr camera_module_cache_reg_ram_181__6 (.Q (camera_module_cache_ram_181__6)
         , .QB (\$dummy [117]), .D (nx18323), .CLK (clk), .R (rst)) ;
    mux21_ni ix18324 (.Y (nx18323), .A0 (camera_module_cache_ram_181__6), .A1 (
             nx35544), .S0 (nx34740)) ;
    dffr camera_module_cache_reg_ram_165__6 (.Q (camera_module_cache_ram_165__6)
         , .QB (\$dummy [118]), .D (nx18333), .CLK (clk), .R (rst)) ;
    mux21_ni ix18334 (.Y (nx18333), .A0 (camera_module_cache_ram_165__6), .A1 (
             nx35546), .S0 (nx34744)) ;
    aoi22 ix23812 (.Y (nx23811), .A0 (camera_module_cache_ram_197__6), .A1 (
          nx36288), .B0 (camera_module_cache_ram_213__6), .B1 (nx36328)) ;
    dffr camera_module_cache_reg_ram_197__6 (.Q (camera_module_cache_ram_197__6)
         , .QB (\$dummy [119]), .D (nx18313), .CLK (clk), .R (rst)) ;
    mux21_ni ix18314 (.Y (nx18313), .A0 (camera_module_cache_ram_197__6), .A1 (
             nx35546), .S0 (nx34736)) ;
    dffr camera_module_cache_reg_ram_213__6 (.Q (camera_module_cache_ram_213__6)
         , .QB (\$dummy [120]), .D (nx18303), .CLK (clk), .R (rst)) ;
    mux21_ni ix18304 (.Y (nx18303), .A0 (camera_module_cache_ram_213__6), .A1 (
             nx35546), .S0 (nx34732)) ;
    aoi22 ix23823 (.Y (nx23822), .A0 (camera_module_cache_ram_229__6), .A1 (
          nx36368), .B0 (camera_module_cache_ram_245__6), .B1 (nx36408)) ;
    dffr camera_module_cache_reg_ram_229__6 (.Q (camera_module_cache_ram_229__6)
         , .QB (\$dummy [121]), .D (nx18293), .CLK (clk), .R (rst)) ;
    mux21_ni ix18294 (.Y (nx18293), .A0 (camera_module_cache_ram_229__6), .A1 (
             nx35546), .S0 (nx34728)) ;
    dffr camera_module_cache_reg_ram_245__6 (.Q (camera_module_cache_ram_245__6)
         , .QB (\$dummy [122]), .D (nx18283), .CLK (clk), .R (rst)) ;
    mux21_ni ix18284 (.Y (nx18283), .A0 (camera_module_cache_ram_245__6), .A1 (
             nx35546), .S0 (nx34724)) ;
    oai21 ix23836 (.Y (nx23835), .A0 (nx21598), .A1 (nx21520), .B0 (nx36472)) ;
    nand04 ix21599 (.Y (nx21598), .A0 (nx23839), .A1 (nx23852), .A2 (nx23863), .A3 (
           nx23875)) ;
    aoi22 ix23840 (.Y (nx23839), .A0 (camera_module_cache_ram_6__6), .A1 (
          nx37030), .B0 (camera_module_cache_ram_22__6), .B1 (nx37032)) ;
    dffr camera_module_cache_reg_ram_6__6 (.Q (camera_module_cache_ram_6__6), .QB (
         \$dummy [123]), .D (nx18273), .CLK (clk), .R (rst)) ;
    mux21_ni ix18274 (.Y (nx18273), .A0 (camera_module_cache_ram_6__6), .A1 (
             nx35546), .S0 (nx34714)) ;
    nand02 ix3889 (.Y (nx3888), .A0 (nx23639), .A1 (nx23423)) ;
    dffr camera_module_cache_reg_ram_22__6 (.Q (camera_module_cache_ram_22__6), 
         .QB (\$dummy [124]), .D (nx18263), .CLK (clk), .R (rst)) ;
    mux21_ni ix18264 (.Y (nx18263), .A0 (camera_module_cache_ram_22__6), .A1 (
             nx35546), .S0 (nx34710)) ;
    aoi22 ix23853 (.Y (nx23852), .A0 (camera_module_cache_ram_38__6), .A1 (
          nx37034), .B0 (camera_module_cache_ram_54__6), .B1 (nx37036)) ;
    dffr camera_module_cache_reg_ram_38__6 (.Q (camera_module_cache_ram_38__6), 
         .QB (\$dummy [125]), .D (nx18253), .CLK (clk), .R (rst)) ;
    mux21_ni ix18254 (.Y (nx18253), .A0 (camera_module_cache_ram_38__6), .A1 (
             nx35548), .S0 (nx34706)) ;
    dffr camera_module_cache_reg_ram_54__6 (.Q (camera_module_cache_ram_54__6), 
         .QB (\$dummy [126]), .D (nx18243), .CLK (clk), .R (rst)) ;
    mux21_ni ix18244 (.Y (nx18243), .A0 (camera_module_cache_ram_54__6), .A1 (
             nx35548), .S0 (nx34702)) ;
    aoi22 ix23864 (.Y (nx23863), .A0 (camera_module_cache_ram_70__6), .A1 (
          nx37038), .B0 (camera_module_cache_ram_86__6), .B1 (nx37040)) ;
    dffr camera_module_cache_reg_ram_70__6 (.Q (camera_module_cache_ram_70__6), 
         .QB (\$dummy [127]), .D (nx18233), .CLK (clk), .R (rst)) ;
    mux21_ni ix18234 (.Y (nx18233), .A0 (camera_module_cache_ram_70__6), .A1 (
             nx35548), .S0 (nx34698)) ;
    dffr camera_module_cache_reg_ram_86__6 (.Q (camera_module_cache_ram_86__6), 
         .QB (\$dummy [128]), .D (nx18223), .CLK (clk), .R (rst)) ;
    mux21_ni ix18224 (.Y (nx18223), .A0 (camera_module_cache_ram_86__6), .A1 (
             nx35548), .S0 (nx34694)) ;
    aoi22 ix23876 (.Y (nx23875), .A0 (camera_module_cache_ram_118__6), .A1 (
          nx37042), .B0 (camera_module_cache_ram_102__6), .B1 (nx37044)) ;
    dffr camera_module_cache_reg_ram_118__6 (.Q (camera_module_cache_ram_118__6)
         , .QB (\$dummy [129]), .D (nx18203), .CLK (clk), .R (rst)) ;
    mux21_ni ix18204 (.Y (nx18203), .A0 (camera_module_cache_ram_118__6), .A1 (
             nx35548), .S0 (nx34686)) ;
    dffr camera_module_cache_reg_ram_102__6 (.Q (camera_module_cache_ram_102__6)
         , .QB (\$dummy [130]), .D (nx18213), .CLK (clk), .R (rst)) ;
    mux21_ni ix18214 (.Y (nx18213), .A0 (camera_module_cache_ram_102__6), .A1 (
             nx35548), .S0 (nx34690)) ;
    nand04 ix21521 (.Y (nx21520), .A0 (nx23889), .A1 (nx23900), .A2 (nx23913), .A3 (
           nx23925)) ;
    aoi22 ix23890 (.Y (nx23889), .A0 (camera_module_cache_ram_134__6), .A1 (
          nx37046), .B0 (camera_module_cache_ram_150__6), .B1 (nx37048)) ;
    dffr camera_module_cache_reg_ram_134__6 (.Q (camera_module_cache_ram_134__6)
         , .QB (\$dummy [131]), .D (nx18193), .CLK (clk), .R (rst)) ;
    mux21_ni ix18194 (.Y (nx18193), .A0 (camera_module_cache_ram_134__6), .A1 (
             nx35548), .S0 (nx34682)) ;
    dffr camera_module_cache_reg_ram_150__6 (.Q (camera_module_cache_ram_150__6)
         , .QB (\$dummy [132]), .D (nx18183), .CLK (clk), .R (rst)) ;
    mux21_ni ix18184 (.Y (nx18183), .A0 (camera_module_cache_ram_150__6), .A1 (
             nx35550), .S0 (nx34678)) ;
    aoi22 ix23901 (.Y (nx23900), .A0 (camera_module_cache_ram_182__6), .A1 (
          nx37050), .B0 (camera_module_cache_ram_166__6), .B1 (nx37052)) ;
    dffr camera_module_cache_reg_ram_182__6 (.Q (camera_module_cache_ram_182__6)
         , .QB (\$dummy [133]), .D (nx18163), .CLK (clk), .R (rst)) ;
    mux21_ni ix18164 (.Y (nx18163), .A0 (camera_module_cache_ram_182__6), .A1 (
             nx35550), .S0 (nx34670)) ;
    dffr camera_module_cache_reg_ram_166__6 (.Q (camera_module_cache_ram_166__6)
         , .QB (\$dummy [134]), .D (nx18173), .CLK (clk), .R (rst)) ;
    mux21_ni ix18174 (.Y (nx18173), .A0 (camera_module_cache_ram_166__6), .A1 (
             nx35550), .S0 (nx34674)) ;
    aoi22 ix23914 (.Y (nx23913), .A0 (camera_module_cache_ram_198__6), .A1 (
          nx36288), .B0 (camera_module_cache_ram_214__6), .B1 (nx36328)) ;
    dffr camera_module_cache_reg_ram_198__6 (.Q (camera_module_cache_ram_198__6)
         , .QB (\$dummy [135]), .D (nx18153), .CLK (clk), .R (rst)) ;
    mux21_ni ix18154 (.Y (nx18153), .A0 (camera_module_cache_ram_198__6), .A1 (
             nx35550), .S0 (nx34666)) ;
    dffr camera_module_cache_reg_ram_214__6 (.Q (camera_module_cache_ram_214__6)
         , .QB (\$dummy [136]), .D (nx18143), .CLK (clk), .R (rst)) ;
    mux21_ni ix18144 (.Y (nx18143), .A0 (camera_module_cache_ram_214__6), .A1 (
             nx35550), .S0 (nx34662)) ;
    aoi22 ix23926 (.Y (nx23925), .A0 (camera_module_cache_ram_230__6), .A1 (
          nx36368), .B0 (camera_module_cache_ram_246__6), .B1 (nx36408)) ;
    dffr camera_module_cache_reg_ram_230__6 (.Q (camera_module_cache_ram_230__6)
         , .QB (\$dummy [137]), .D (nx18133), .CLK (clk), .R (rst)) ;
    mux21_ni ix18134 (.Y (nx18133), .A0 (camera_module_cache_ram_230__6), .A1 (
             nx35550), .S0 (nx34658)) ;
    dffr camera_module_cache_reg_ram_246__6 (.Q (camera_module_cache_ram_246__6)
         , .QB (\$dummy [138]), .D (nx18123), .CLK (clk), .R (rst)) ;
    mux21_ni ix18124 (.Y (nx18123), .A0 (camera_module_cache_ram_246__6), .A1 (
             nx35550), .S0 (nx34654)) ;
    oai21 ix23939 (.Y (nx23938), .A0 (nx21436), .A1 (nx21358), .B0 (nx36476)) ;
    nand04 ix21437 (.Y (nx21436), .A0 (nx23941), .A1 (nx23954), .A2 (nx23966), .A3 (
           nx23977)) ;
    aoi22 ix23942 (.Y (nx23941), .A0 (camera_module_cache_ram_7__6), .A1 (
          nx35810), .B0 (camera_module_cache_ram_23__6), .B1 (nx35850)) ;
    dffr camera_module_cache_reg_ram_7__6 (.Q (camera_module_cache_ram_7__6), .QB (
         \$dummy [139]), .D (nx18113), .CLK (clk), .R (rst)) ;
    mux21_ni ix18114 (.Y (nx18113), .A0 (camera_module_cache_ram_7__6), .A1 (
             nx35552), .S0 (nx34644)) ;
    nand02 ix3597 (.Y (nx3596), .A0 (nx23639), .A1 (nx23529)) ;
    dffr camera_module_cache_reg_ram_23__6 (.Q (camera_module_cache_ram_23__6), 
         .QB (\$dummy [140]), .D (nx18103), .CLK (clk), .R (rst)) ;
    mux21_ni ix18104 (.Y (nx18103), .A0 (camera_module_cache_ram_23__6), .A1 (
             nx35552), .S0 (nx34640)) ;
    aoi22 ix23955 (.Y (nx23954), .A0 (camera_module_cache_ram_39__6), .A1 (
          nx35890), .B0 (camera_module_cache_ram_55__6), .B1 (nx35930)) ;
    dffr camera_module_cache_reg_ram_39__6 (.Q (camera_module_cache_ram_39__6), 
         .QB (\$dummy [141]), .D (nx18093), .CLK (clk), .R (rst)) ;
    mux21_ni ix18094 (.Y (nx18093), .A0 (camera_module_cache_ram_39__6), .A1 (
             nx35552), .S0 (nx34636)) ;
    dffr camera_module_cache_reg_ram_55__6 (.Q (camera_module_cache_ram_55__6), 
         .QB (\$dummy [142]), .D (nx18083), .CLK (clk), .R (rst)) ;
    mux21_ni ix18084 (.Y (nx18083), .A0 (camera_module_cache_ram_55__6), .A1 (
             nx35552), .S0 (nx34632)) ;
    aoi22 ix23967 (.Y (nx23966), .A0 (camera_module_cache_ram_71__6), .A1 (
          nx35970), .B0 (camera_module_cache_ram_87__6), .B1 (nx36010)) ;
    dffr camera_module_cache_reg_ram_71__6 (.Q (camera_module_cache_ram_71__6), 
         .QB (\$dummy [143]), .D (nx18073), .CLK (clk), .R (rst)) ;
    mux21_ni ix18074 (.Y (nx18073), .A0 (camera_module_cache_ram_71__6), .A1 (
             nx35552), .S0 (nx34628)) ;
    dffr camera_module_cache_reg_ram_87__6 (.Q (camera_module_cache_ram_87__6), 
         .QB (\$dummy [144]), .D (nx18063), .CLK (clk), .R (rst)) ;
    mux21_ni ix18064 (.Y (nx18063), .A0 (camera_module_cache_ram_87__6), .A1 (
             nx35552), .S0 (nx34624)) ;
    aoi22 ix23978 (.Y (nx23977), .A0 (camera_module_cache_ram_119__6), .A1 (
          nx36050), .B0 (camera_module_cache_ram_103__6), .B1 (nx36090)) ;
    dffr camera_module_cache_reg_ram_119__6 (.Q (camera_module_cache_ram_119__6)
         , .QB (\$dummy [145]), .D (nx18043), .CLK (clk), .R (rst)) ;
    mux21_ni ix18044 (.Y (nx18043), .A0 (camera_module_cache_ram_119__6), .A1 (
             nx35552), .S0 (nx34616)) ;
    dffr camera_module_cache_reg_ram_103__6 (.Q (camera_module_cache_ram_103__6)
         , .QB (\$dummy [146]), .D (nx18053), .CLK (clk), .R (rst)) ;
    mux21_ni ix18054 (.Y (nx18053), .A0 (camera_module_cache_ram_103__6), .A1 (
             nx35554), .S0 (nx34620)) ;
    nand04 ix21359 (.Y (nx21358), .A0 (nx23989), .A1 (nx24001), .A2 (nx24012), .A3 (
           nx24024)) ;
    aoi22 ix23990 (.Y (nx23989), .A0 (camera_module_cache_ram_135__6), .A1 (
          nx36130), .B0 (camera_module_cache_ram_151__6), .B1 (nx36170)) ;
    dffr camera_module_cache_reg_ram_135__6 (.Q (camera_module_cache_ram_135__6)
         , .QB (\$dummy [147]), .D (nx18033), .CLK (clk), .R (rst)) ;
    mux21_ni ix18034 (.Y (nx18033), .A0 (camera_module_cache_ram_135__6), .A1 (
             nx35554), .S0 (nx34612)) ;
    dffr camera_module_cache_reg_ram_151__6 (.Q (camera_module_cache_ram_151__6)
         , .QB (\$dummy [148]), .D (nx18023), .CLK (clk), .R (rst)) ;
    mux21_ni ix18024 (.Y (nx18023), .A0 (camera_module_cache_ram_151__6), .A1 (
             nx35554), .S0 (nx34608)) ;
    aoi22 ix24002 (.Y (nx24001), .A0 (camera_module_cache_ram_183__6), .A1 (
          nx36210), .B0 (camera_module_cache_ram_167__6), .B1 (nx36250)) ;
    dffr camera_module_cache_reg_ram_183__6 (.Q (camera_module_cache_ram_183__6)
         , .QB (\$dummy [149]), .D (nx18003), .CLK (clk), .R (rst)) ;
    mux21_ni ix18004 (.Y (nx18003), .A0 (camera_module_cache_ram_183__6), .A1 (
             nx35554), .S0 (nx34600)) ;
    dffr camera_module_cache_reg_ram_167__6 (.Q (camera_module_cache_ram_167__6)
         , .QB (\$dummy [150]), .D (nx18013), .CLK (clk), .R (rst)) ;
    mux21_ni ix18014 (.Y (nx18013), .A0 (camera_module_cache_ram_167__6), .A1 (
             nx35554), .S0 (nx34604)) ;
    aoi22 ix24013 (.Y (nx24012), .A0 (camera_module_cache_ram_199__6), .A1 (
          nx36290), .B0 (camera_module_cache_ram_215__6), .B1 (nx36330)) ;
    dffr camera_module_cache_reg_ram_199__6 (.Q (camera_module_cache_ram_199__6)
         , .QB (\$dummy [151]), .D (nx17993), .CLK (clk), .R (rst)) ;
    mux21_ni ix17994 (.Y (nx17993), .A0 (camera_module_cache_ram_199__6), .A1 (
             nx35554), .S0 (nx34596)) ;
    dffr camera_module_cache_reg_ram_215__6 (.Q (camera_module_cache_ram_215__6)
         , .QB (\$dummy [152]), .D (nx17983), .CLK (clk), .R (rst)) ;
    mux21_ni ix17984 (.Y (nx17983), .A0 (camera_module_cache_ram_215__6), .A1 (
             nx35554), .S0 (nx34592)) ;
    aoi22 ix24025 (.Y (nx24024), .A0 (camera_module_cache_ram_231__6), .A1 (
          nx36370), .B0 (camera_module_cache_ram_247__6), .B1 (nx36410)) ;
    dffr camera_module_cache_reg_ram_231__6 (.Q (camera_module_cache_ram_231__6)
         , .QB (\$dummy [153]), .D (nx17973), .CLK (clk), .R (rst)) ;
    mux21_ni ix17974 (.Y (nx17973), .A0 (camera_module_cache_ram_231__6), .A1 (
             nx35556), .S0 (nx34588)) ;
    dffr camera_module_cache_reg_ram_247__6 (.Q (camera_module_cache_ram_247__6)
         , .QB (\$dummy [154]), .D (nx17963), .CLK (clk), .R (rst)) ;
    mux21_ni ix17964 (.Y (nx17963), .A0 (camera_module_cache_ram_247__6), .A1 (
             nx35556), .S0 (nx34584)) ;
    nand04 ix21279 (.Y (nx21278), .A0 (nx24041), .A1 (nx24146), .A2 (nx24248), .A3 (
           nx24349)) ;
    oai21 ix24042 (.Y (nx24041), .A0 (nx21268), .A1 (nx21190), .B0 (nx36480)) ;
    nand04 ix21269 (.Y (nx21268), .A0 (nx24045), .A1 (nx24060), .A2 (nx24073), .A3 (
           nx24084)) ;
    aoi22 ix24046 (.Y (nx24045), .A0 (camera_module_cache_ram_8__6), .A1 (
          nx35810), .B0 (camera_module_cache_ram_24__6), .B1 (nx35850)) ;
    dffr camera_module_cache_reg_ram_8__6 (.Q (camera_module_cache_ram_8__6), .QB (
         \$dummy [155]), .D (nx17953), .CLK (clk), .R (rst)) ;
    mux21_ni ix17954 (.Y (nx17953), .A0 (camera_module_cache_ram_8__6), .A1 (
             nx35556), .S0 (nx34574)) ;
    nand02 ix3295 (.Y (nx3294), .A0 (nx24053), .A1 (nx23105)) ;
    dffr camera_module_cache_reg_ram_24__6 (.Q (camera_module_cache_ram_24__6), 
         .QB (\$dummy [156]), .D (nx17943), .CLK (clk), .R (rst)) ;
    mux21_ni ix17944 (.Y (nx17943), .A0 (camera_module_cache_ram_24__6), .A1 (
             nx35556), .S0 (nx34570)) ;
    aoi22 ix24061 (.Y (nx24060), .A0 (camera_module_cache_ram_40__6), .A1 (
          nx35890), .B0 (camera_module_cache_ram_56__6), .B1 (nx35930)) ;
    dffr camera_module_cache_reg_ram_40__6 (.Q (camera_module_cache_ram_40__6), 
         .QB (\$dummy [157]), .D (nx17933), .CLK (clk), .R (rst)) ;
    mux21_ni ix17934 (.Y (nx17933), .A0 (camera_module_cache_ram_40__6), .A1 (
             nx35556), .S0 (nx34566)) ;
    dffr camera_module_cache_reg_ram_56__6 (.Q (camera_module_cache_ram_56__6), 
         .QB (\$dummy [158]), .D (nx17923), .CLK (clk), .R (rst)) ;
    mux21_ni ix17924 (.Y (nx17923), .A0 (camera_module_cache_ram_56__6), .A1 (
             nx35556), .S0 (nx34562)) ;
    aoi22 ix24074 (.Y (nx24073), .A0 (camera_module_cache_ram_72__6), .A1 (
          nx35970), .B0 (camera_module_cache_ram_88__6), .B1 (nx36010)) ;
    dffr camera_module_cache_reg_ram_72__6 (.Q (camera_module_cache_ram_72__6), 
         .QB (\$dummy [159]), .D (nx17913), .CLK (clk), .R (rst)) ;
    mux21_ni ix17914 (.Y (nx17913), .A0 (camera_module_cache_ram_72__6), .A1 (
             nx35556), .S0 (nx34558)) ;
    dffr camera_module_cache_reg_ram_88__6 (.Q (camera_module_cache_ram_88__6), 
         .QB (\$dummy [160]), .D (nx17903), .CLK (clk), .R (rst)) ;
    mux21_ni ix17904 (.Y (nx17903), .A0 (camera_module_cache_ram_88__6), .A1 (
             nx35558), .S0 (nx34554)) ;
    aoi22 ix24085 (.Y (nx24084), .A0 (camera_module_cache_ram_120__6), .A1 (
          nx36050), .B0 (camera_module_cache_ram_104__6), .B1 (nx36090)) ;
    dffr camera_module_cache_reg_ram_120__6 (.Q (camera_module_cache_ram_120__6)
         , .QB (\$dummy [161]), .D (nx17883), .CLK (clk), .R (rst)) ;
    mux21_ni ix17884 (.Y (nx17883), .A0 (camera_module_cache_ram_120__6), .A1 (
             nx35558), .S0 (nx34546)) ;
    dffr camera_module_cache_reg_ram_104__6 (.Q (camera_module_cache_ram_104__6)
         , .QB (\$dummy [162]), .D (nx17893), .CLK (clk), .R (rst)) ;
    mux21_ni ix17894 (.Y (nx17893), .A0 (camera_module_cache_ram_104__6), .A1 (
             nx35558), .S0 (nx34550)) ;
    nand04 ix21191 (.Y (nx21190), .A0 (nx24097), .A1 (nx24109), .A2 (nx24120), .A3 (
           nx24133)) ;
    aoi22 ix24098 (.Y (nx24097), .A0 (camera_module_cache_ram_136__6), .A1 (
          nx36130), .B0 (camera_module_cache_ram_152__6), .B1 (nx36170)) ;
    dffr camera_module_cache_reg_ram_136__6 (.Q (camera_module_cache_ram_136__6)
         , .QB (\$dummy [163]), .D (nx17873), .CLK (clk), .R (rst)) ;
    mux21_ni ix17874 (.Y (nx17873), .A0 (camera_module_cache_ram_136__6), .A1 (
             nx35558), .S0 (nx34542)) ;
    dffr camera_module_cache_reg_ram_152__6 (.Q (camera_module_cache_ram_152__6)
         , .QB (\$dummy [164]), .D (nx17863), .CLK (clk), .R (rst)) ;
    mux21_ni ix17864 (.Y (nx17863), .A0 (camera_module_cache_ram_152__6), .A1 (
             nx35558), .S0 (nx34538)) ;
    aoi22 ix24110 (.Y (nx24109), .A0 (camera_module_cache_ram_184__6), .A1 (
          nx36210), .B0 (camera_module_cache_ram_168__6), .B1 (nx36250)) ;
    dffr camera_module_cache_reg_ram_184__6 (.Q (camera_module_cache_ram_184__6)
         , .QB (\$dummy [165]), .D (nx17843), .CLK (clk), .R (rst)) ;
    mux21_ni ix17844 (.Y (nx17843), .A0 (camera_module_cache_ram_184__6), .A1 (
             nx35558), .S0 (nx34530)) ;
    dffr camera_module_cache_reg_ram_168__6 (.Q (camera_module_cache_ram_168__6)
         , .QB (\$dummy [166]), .D (nx17853), .CLK (clk), .R (rst)) ;
    mux21_ni ix17854 (.Y (nx17853), .A0 (camera_module_cache_ram_168__6), .A1 (
             nx35558), .S0 (nx34534)) ;
    aoi22 ix24121 (.Y (nx24120), .A0 (camera_module_cache_ram_200__6), .A1 (
          nx36290), .B0 (camera_module_cache_ram_216__6), .B1 (nx36330)) ;
    dffr camera_module_cache_reg_ram_200__6 (.Q (camera_module_cache_ram_200__6)
         , .QB (\$dummy [167]), .D (nx17833), .CLK (clk), .R (rst)) ;
    mux21_ni ix17834 (.Y (nx17833), .A0 (camera_module_cache_ram_200__6), .A1 (
             nx35560), .S0 (nx34526)) ;
    dffr camera_module_cache_reg_ram_216__6 (.Q (camera_module_cache_ram_216__6)
         , .QB (\$dummy [168]), .D (nx17823), .CLK (clk), .R (rst)) ;
    mux21_ni ix17824 (.Y (nx17823), .A0 (camera_module_cache_ram_216__6), .A1 (
             nx35560), .S0 (nx34522)) ;
    aoi22 ix24134 (.Y (nx24133), .A0 (camera_module_cache_ram_232__6), .A1 (
          nx36370), .B0 (camera_module_cache_ram_248__6), .B1 (nx36410)) ;
    dffr camera_module_cache_reg_ram_232__6 (.Q (camera_module_cache_ram_232__6)
         , .QB (\$dummy [169]), .D (nx17813), .CLK (clk), .R (rst)) ;
    mux21_ni ix17814 (.Y (nx17813), .A0 (camera_module_cache_ram_232__6), .A1 (
             nx35560), .S0 (nx34518)) ;
    dffr camera_module_cache_reg_ram_248__6 (.Q (camera_module_cache_ram_248__6)
         , .QB (\$dummy [170]), .D (nx17803), .CLK (clk), .R (rst)) ;
    mux21_ni ix17804 (.Y (nx17803), .A0 (camera_module_cache_ram_248__6), .A1 (
             nx35560), .S0 (nx34514)) ;
    oai21 ix24147 (.Y (nx24146), .A0 (nx21106), .A1 (nx21028), .B0 (nx36484)) ;
    nand04 ix21107 (.Y (nx21106), .A0 (nx24149), .A1 (nx24162), .A2 (nx24174), .A3 (
           nx24184)) ;
    aoi22 ix24150 (.Y (nx24149), .A0 (camera_module_cache_ram_9__6), .A1 (
          nx35810), .B0 (camera_module_cache_ram_25__6), .B1 (nx35850)) ;
    dffr camera_module_cache_reg_ram_9__6 (.Q (camera_module_cache_ram_9__6), .QB (
         \$dummy [171]), .D (nx17793), .CLK (clk), .R (rst)) ;
    mux21_ni ix17794 (.Y (nx17793), .A0 (camera_module_cache_ram_9__6), .A1 (
             nx35560), .S0 (nx34504)) ;
    nand02 ix3003 (.Y (nx3002), .A0 (nx24053), .A1 (nx23314)) ;
    dffr camera_module_cache_reg_ram_25__6 (.Q (camera_module_cache_ram_25__6), 
         .QB (\$dummy [172]), .D (nx17783), .CLK (clk), .R (rst)) ;
    mux21_ni ix17784 (.Y (nx17783), .A0 (camera_module_cache_ram_25__6), .A1 (
             nx35560), .S0 (nx34500)) ;
    aoi22 ix24163 (.Y (nx24162), .A0 (camera_module_cache_ram_41__6), .A1 (
          nx35890), .B0 (camera_module_cache_ram_57__6), .B1 (nx35930)) ;
    dffr camera_module_cache_reg_ram_41__6 (.Q (camera_module_cache_ram_41__6), 
         .QB (\$dummy [173]), .D (nx17773), .CLK (clk), .R (rst)) ;
    mux21_ni ix17774 (.Y (nx17773), .A0 (camera_module_cache_ram_41__6), .A1 (
             nx35560), .S0 (nx34496)) ;
    dffr camera_module_cache_reg_ram_57__6 (.Q (camera_module_cache_ram_57__6), 
         .QB (\$dummy [174]), .D (nx17763), .CLK (clk), .R (rst)) ;
    mux21_ni ix17764 (.Y (nx17763), .A0 (camera_module_cache_ram_57__6), .A1 (
             nx35562), .S0 (nx34492)) ;
    aoi22 ix24175 (.Y (nx24174), .A0 (camera_module_cache_ram_73__6), .A1 (
          nx35970), .B0 (camera_module_cache_ram_89__6), .B1 (nx36010)) ;
    dffr camera_module_cache_reg_ram_73__6 (.Q (camera_module_cache_ram_73__6), 
         .QB (\$dummy [175]), .D (nx17753), .CLK (clk), .R (rst)) ;
    mux21_ni ix17754 (.Y (nx17753), .A0 (camera_module_cache_ram_73__6), .A1 (
             nx35562), .S0 (nx34488)) ;
    dffr camera_module_cache_reg_ram_89__6 (.Q (camera_module_cache_ram_89__6), 
         .QB (\$dummy [176]), .D (nx17743), .CLK (clk), .R (rst)) ;
    mux21_ni ix17744 (.Y (nx17743), .A0 (camera_module_cache_ram_89__6), .A1 (
             nx35562), .S0 (nx34484)) ;
    aoi22 ix24185 (.Y (nx24184), .A0 (camera_module_cache_ram_121__6), .A1 (
          nx36050), .B0 (camera_module_cache_ram_105__6), .B1 (nx36090)) ;
    dffr camera_module_cache_reg_ram_121__6 (.Q (camera_module_cache_ram_121__6)
         , .QB (\$dummy [177]), .D (nx17723), .CLK (clk), .R (rst)) ;
    mux21_ni ix17724 (.Y (nx17723), .A0 (camera_module_cache_ram_121__6), .A1 (
             nx35562), .S0 (nx34476)) ;
    dffr camera_module_cache_reg_ram_105__6 (.Q (camera_module_cache_ram_105__6)
         , .QB (\$dummy [178]), .D (nx17733), .CLK (clk), .R (rst)) ;
    mux21_ni ix17734 (.Y (nx17733), .A0 (camera_module_cache_ram_105__6), .A1 (
             nx35562), .S0 (nx34480)) ;
    nand04 ix21029 (.Y (nx21028), .A0 (nx24197), .A1 (nx24209), .A2 (nx24222), .A3 (
           nx24235)) ;
    aoi22 ix24198 (.Y (nx24197), .A0 (camera_module_cache_ram_137__6), .A1 (
          nx36130), .B0 (camera_module_cache_ram_153__6), .B1 (nx36170)) ;
    dffr camera_module_cache_reg_ram_137__6 (.Q (camera_module_cache_ram_137__6)
         , .QB (\$dummy [179]), .D (nx17713), .CLK (clk), .R (rst)) ;
    mux21_ni ix17714 (.Y (nx17713), .A0 (camera_module_cache_ram_137__6), .A1 (
             nx35562), .S0 (nx34472)) ;
    dffr camera_module_cache_reg_ram_153__6 (.Q (camera_module_cache_ram_153__6)
         , .QB (\$dummy [180]), .D (nx17703), .CLK (clk), .R (rst)) ;
    mux21_ni ix17704 (.Y (nx17703), .A0 (camera_module_cache_ram_153__6), .A1 (
             nx35562), .S0 (nx34468)) ;
    aoi22 ix24210 (.Y (nx24209), .A0 (camera_module_cache_ram_185__6), .A1 (
          nx36210), .B0 (camera_module_cache_ram_169__6), .B1 (nx36250)) ;
    dffr camera_module_cache_reg_ram_185__6 (.Q (camera_module_cache_ram_185__6)
         , .QB (\$dummy [181]), .D (nx17683), .CLK (clk), .R (rst)) ;
    mux21_ni ix17684 (.Y (nx17683), .A0 (camera_module_cache_ram_185__6), .A1 (
             nx35564), .S0 (nx34460)) ;
    dffr camera_module_cache_reg_ram_169__6 (.Q (camera_module_cache_ram_169__6)
         , .QB (\$dummy [182]), .D (nx17693), .CLK (clk), .R (rst)) ;
    mux21_ni ix17694 (.Y (nx17693), .A0 (camera_module_cache_ram_169__6), .A1 (
             nx35564), .S0 (nx34464)) ;
    aoi22 ix24223 (.Y (nx24222), .A0 (camera_module_cache_ram_201__6), .A1 (
          nx36290), .B0 (camera_module_cache_ram_217__6), .B1 (nx36330)) ;
    dffr camera_module_cache_reg_ram_201__6 (.Q (camera_module_cache_ram_201__6)
         , .QB (\$dummy [183]), .D (nx17673), .CLK (clk), .R (rst)) ;
    mux21_ni ix17674 (.Y (nx17673), .A0 (camera_module_cache_ram_201__6), .A1 (
             nx35564), .S0 (nx34456)) ;
    dffr camera_module_cache_reg_ram_217__6 (.Q (camera_module_cache_ram_217__6)
         , .QB (\$dummy [184]), .D (nx17663), .CLK (clk), .R (rst)) ;
    mux21_ni ix17664 (.Y (nx17663), .A0 (camera_module_cache_ram_217__6), .A1 (
             nx35564), .S0 (nx34452)) ;
    aoi22 ix24236 (.Y (nx24235), .A0 (camera_module_cache_ram_233__6), .A1 (
          nx36370), .B0 (camera_module_cache_ram_249__6), .B1 (nx36410)) ;
    dffr camera_module_cache_reg_ram_233__6 (.Q (camera_module_cache_ram_233__6)
         , .QB (\$dummy [185]), .D (nx17653), .CLK (clk), .R (rst)) ;
    mux21_ni ix17654 (.Y (nx17653), .A0 (camera_module_cache_ram_233__6), .A1 (
             nx35564), .S0 (nx34448)) ;
    dffr camera_module_cache_reg_ram_249__6 (.Q (camera_module_cache_ram_249__6)
         , .QB (\$dummy [186]), .D (nx17643), .CLK (clk), .R (rst)) ;
    mux21_ni ix17644 (.Y (nx17643), .A0 (camera_module_cache_ram_249__6), .A1 (
             nx35564), .S0 (nx34444)) ;
    oai21 ix24249 (.Y (nx24248), .A0 (nx20942), .A1 (nx20864), .B0 (nx36488)) ;
    nand04 ix20943 (.Y (nx20942), .A0 (nx24251), .A1 (nx24264), .A2 (nx24276), .A3 (
           nx24286)) ;
    aoi22 ix24252 (.Y (nx24251), .A0 (camera_module_cache_ram_10__6), .A1 (
          nx35810), .B0 (camera_module_cache_ram_26__6), .B1 (nx35850)) ;
    dffr camera_module_cache_reg_ram_10__6 (.Q (camera_module_cache_ram_10__6), 
         .QB (\$dummy [187]), .D (nx17633), .CLK (clk), .R (rst)) ;
    mux21_ni ix17634 (.Y (nx17633), .A0 (camera_module_cache_ram_10__6), .A1 (
             nx35564), .S0 (nx34434)) ;
    nand02 ix2709 (.Y (nx2708), .A0 (nx24053), .A1 (nx23423)) ;
    dffr camera_module_cache_reg_ram_26__6 (.Q (camera_module_cache_ram_26__6), 
         .QB (\$dummy [188]), .D (nx17623), .CLK (clk), .R (rst)) ;
    mux21_ni ix17624 (.Y (nx17623), .A0 (camera_module_cache_ram_26__6), .A1 (
             nx35566), .S0 (nx34430)) ;
    aoi22 ix24265 (.Y (nx24264), .A0 (camera_module_cache_ram_42__6), .A1 (
          nx35890), .B0 (camera_module_cache_ram_58__6), .B1 (nx35930)) ;
    dffr camera_module_cache_reg_ram_42__6 (.Q (camera_module_cache_ram_42__6), 
         .QB (\$dummy [189]), .D (nx17613), .CLK (clk), .R (rst)) ;
    mux21_ni ix17614 (.Y (nx17613), .A0 (camera_module_cache_ram_42__6), .A1 (
             nx35566), .S0 (nx34426)) ;
    dffr camera_module_cache_reg_ram_58__6 (.Q (camera_module_cache_ram_58__6), 
         .QB (\$dummy [190]), .D (nx17603), .CLK (clk), .R (rst)) ;
    mux21_ni ix17604 (.Y (nx17603), .A0 (camera_module_cache_ram_58__6), .A1 (
             nx35566), .S0 (nx34422)) ;
    aoi22 ix24277 (.Y (nx24276), .A0 (camera_module_cache_ram_74__6), .A1 (
          nx35970), .B0 (camera_module_cache_ram_90__6), .B1 (nx36010)) ;
    dffr camera_module_cache_reg_ram_74__6 (.Q (camera_module_cache_ram_74__6), 
         .QB (\$dummy [191]), .D (nx17593), .CLK (clk), .R (rst)) ;
    mux21_ni ix17594 (.Y (nx17593), .A0 (camera_module_cache_ram_74__6), .A1 (
             nx35566), .S0 (nx34418)) ;
    dffr camera_module_cache_reg_ram_90__6 (.Q (camera_module_cache_ram_90__6), 
         .QB (\$dummy [192]), .D (nx17583), .CLK (clk), .R (rst)) ;
    mux21_ni ix17584 (.Y (nx17583), .A0 (camera_module_cache_ram_90__6), .A1 (
             nx35566), .S0 (nx34414)) ;
    aoi22 ix24287 (.Y (nx24286), .A0 (camera_module_cache_ram_122__6), .A1 (
          nx36050), .B0 (camera_module_cache_ram_106__6), .B1 (nx36090)) ;
    dffr camera_module_cache_reg_ram_122__6 (.Q (camera_module_cache_ram_122__6)
         , .QB (\$dummy [193]), .D (nx17563), .CLK (clk), .R (rst)) ;
    mux21_ni ix17564 (.Y (nx17563), .A0 (camera_module_cache_ram_122__6), .A1 (
             nx35566), .S0 (nx34406)) ;
    dffr camera_module_cache_reg_ram_106__6 (.Q (camera_module_cache_ram_106__6)
         , .QB (\$dummy [194]), .D (nx17573), .CLK (clk), .R (rst)) ;
    mux21_ni ix17574 (.Y (nx17573), .A0 (camera_module_cache_ram_106__6), .A1 (
             nx35566), .S0 (nx34410)) ;
    nand04 ix20865 (.Y (nx20864), .A0 (nx24300), .A1 (nx24313), .A2 (nx24324), .A3 (
           nx24336)) ;
    aoi22 ix24301 (.Y (nx24300), .A0 (camera_module_cache_ram_138__6), .A1 (
          nx36130), .B0 (camera_module_cache_ram_154__6), .B1 (nx36170)) ;
    dffr camera_module_cache_reg_ram_138__6 (.Q (camera_module_cache_ram_138__6)
         , .QB (\$dummy [195]), .D (nx17553), .CLK (clk), .R (rst)) ;
    mux21_ni ix17554 (.Y (nx17553), .A0 (camera_module_cache_ram_138__6), .A1 (
             nx35568), .S0 (nx34402)) ;
    dffr camera_module_cache_reg_ram_154__6 (.Q (camera_module_cache_ram_154__6)
         , .QB (\$dummy [196]), .D (nx17543), .CLK (clk), .R (rst)) ;
    mux21_ni ix17544 (.Y (nx17543), .A0 (camera_module_cache_ram_154__6), .A1 (
             nx35568), .S0 (nx34398)) ;
    aoi22 ix24314 (.Y (nx24313), .A0 (camera_module_cache_ram_186__6), .A1 (
          nx36210), .B0 (camera_module_cache_ram_170__6), .B1 (nx36250)) ;
    dffr camera_module_cache_reg_ram_186__6 (.Q (camera_module_cache_ram_186__6)
         , .QB (\$dummy [197]), .D (nx17523), .CLK (clk), .R (rst)) ;
    mux21_ni ix17524 (.Y (nx17523), .A0 (camera_module_cache_ram_186__6), .A1 (
             nx35568), .S0 (nx34390)) ;
    dffr camera_module_cache_reg_ram_170__6 (.Q (camera_module_cache_ram_170__6)
         , .QB (\$dummy [198]), .D (nx17533), .CLK (clk), .R (rst)) ;
    mux21_ni ix17534 (.Y (nx17533), .A0 (camera_module_cache_ram_170__6), .A1 (
             nx35568), .S0 (nx34394)) ;
    aoi22 ix24325 (.Y (nx24324), .A0 (camera_module_cache_ram_202__6), .A1 (
          nx36290), .B0 (camera_module_cache_ram_218__6), .B1 (nx36330)) ;
    dffr camera_module_cache_reg_ram_202__6 (.Q (camera_module_cache_ram_202__6)
         , .QB (\$dummy [199]), .D (nx17513), .CLK (clk), .R (rst)) ;
    mux21_ni ix17514 (.Y (nx17513), .A0 (camera_module_cache_ram_202__6), .A1 (
             nx35568), .S0 (nx34386)) ;
    dffr camera_module_cache_reg_ram_218__6 (.Q (camera_module_cache_ram_218__6)
         , .QB (\$dummy [200]), .D (nx17503), .CLK (clk), .R (rst)) ;
    mux21_ni ix17504 (.Y (nx17503), .A0 (camera_module_cache_ram_218__6), .A1 (
             nx35568), .S0 (nx34382)) ;
    aoi22 ix24337 (.Y (nx24336), .A0 (camera_module_cache_ram_234__6), .A1 (
          nx36370), .B0 (camera_module_cache_ram_250__6), .B1 (nx36410)) ;
    dffr camera_module_cache_reg_ram_234__6 (.Q (camera_module_cache_ram_234__6)
         , .QB (\$dummy [201]), .D (nx17493), .CLK (clk), .R (rst)) ;
    mux21_ni ix17494 (.Y (nx17493), .A0 (camera_module_cache_ram_234__6), .A1 (
             nx35568), .S0 (nx34378)) ;
    dffr camera_module_cache_reg_ram_250__6 (.Q (camera_module_cache_ram_250__6)
         , .QB (\$dummy [202]), .D (nx17483), .CLK (clk), .R (rst)) ;
    mux21_ni ix17484 (.Y (nx17483), .A0 (camera_module_cache_ram_250__6), .A1 (
             nx35570), .S0 (nx34374)) ;
    oai21 ix24350 (.Y (nx24349), .A0 (nx20780), .A1 (nx20702), .B0 (nx36492)) ;
    nand04 ix20781 (.Y (nx20780), .A0 (nx24353), .A1 (nx24364), .A2 (nx24379), .A3 (
           nx24390)) ;
    aoi22 ix24354 (.Y (nx24353), .A0 (camera_module_cache_ram_11__6), .A1 (
          nx35810), .B0 (camera_module_cache_ram_27__6), .B1 (nx35850)) ;
    dffr camera_module_cache_reg_ram_11__6 (.Q (camera_module_cache_ram_11__6), 
         .QB (\$dummy [203]), .D (nx17473), .CLK (clk), .R (rst)) ;
    mux21_ni ix17474 (.Y (nx17473), .A0 (camera_module_cache_ram_11__6), .A1 (
             nx35570), .S0 (nx34364)) ;
    nand02 ix2417 (.Y (nx2416), .A0 (nx24053), .A1 (nx23529)) ;
    dffr camera_module_cache_reg_ram_27__6 (.Q (camera_module_cache_ram_27__6), 
         .QB (\$dummy [204]), .D (nx17463), .CLK (clk), .R (rst)) ;
    mux21_ni ix17464 (.Y (nx17463), .A0 (camera_module_cache_ram_27__6), .A1 (
             nx35570), .S0 (nx34360)) ;
    aoi22 ix24365 (.Y (nx24364), .A0 (camera_module_cache_ram_43__6), .A1 (
          nx35890), .B0 (camera_module_cache_ram_59__6), .B1 (nx35930)) ;
    dffr camera_module_cache_reg_ram_43__6 (.Q (camera_module_cache_ram_43__6), 
         .QB (\$dummy [205]), .D (nx17453), .CLK (clk), .R (rst)) ;
    mux21_ni ix17454 (.Y (nx17453), .A0 (camera_module_cache_ram_43__6), .A1 (
             nx35570), .S0 (nx34356)) ;
    dffr camera_module_cache_reg_ram_59__6 (.Q (camera_module_cache_ram_59__6), 
         .QB (\$dummy [206]), .D (nx17443), .CLK (clk), .R (rst)) ;
    mux21_ni ix17444 (.Y (nx17443), .A0 (camera_module_cache_ram_59__6), .A1 (
             nx35570), .S0 (nx34352)) ;
    aoi22 ix24380 (.Y (nx24379), .A0 (camera_module_cache_ram_75__6), .A1 (
          nx35970), .B0 (camera_module_cache_ram_91__6), .B1 (nx36010)) ;
    dffr camera_module_cache_reg_ram_75__6 (.Q (camera_module_cache_ram_75__6), 
         .QB (\$dummy [207]), .D (nx17433), .CLK (clk), .R (rst)) ;
    mux21_ni ix17434 (.Y (nx17433), .A0 (camera_module_cache_ram_75__6), .A1 (
             nx35570), .S0 (nx34348)) ;
    dffr camera_module_cache_reg_ram_91__6 (.Q (camera_module_cache_ram_91__6), 
         .QB (\$dummy [208]), .D (nx17423), .CLK (clk), .R (rst)) ;
    mux21_ni ix17424 (.Y (nx17423), .A0 (camera_module_cache_ram_91__6), .A1 (
             nx35570), .S0 (nx34344)) ;
    aoi22 ix24391 (.Y (nx24390), .A0 (camera_module_cache_ram_123__6), .A1 (
          nx36050), .B0 (camera_module_cache_ram_107__6), .B1 (nx36090)) ;
    dffr camera_module_cache_reg_ram_123__6 (.Q (camera_module_cache_ram_123__6)
         , .QB (\$dummy [209]), .D (nx17403), .CLK (clk), .R (rst)) ;
    mux21_ni ix17404 (.Y (nx17403), .A0 (camera_module_cache_ram_123__6), .A1 (
             nx35572), .S0 (nx34336)) ;
    dffr camera_module_cache_reg_ram_107__6 (.Q (camera_module_cache_ram_107__6)
         , .QB (\$dummy [210]), .D (nx17413), .CLK (clk), .R (rst)) ;
    mux21_ni ix17414 (.Y (nx17413), .A0 (camera_module_cache_ram_107__6), .A1 (
             nx35572), .S0 (nx34340)) ;
    nand04 ix20703 (.Y (nx20702), .A0 (nx24403), .A1 (nx24415), .A2 (nx24428), .A3 (
           nx24440)) ;
    aoi22 ix24404 (.Y (nx24403), .A0 (camera_module_cache_ram_139__6), .A1 (
          nx36130), .B0 (camera_module_cache_ram_155__6), .B1 (nx36170)) ;
    dffr camera_module_cache_reg_ram_139__6 (.Q (camera_module_cache_ram_139__6)
         , .QB (\$dummy [211]), .D (nx17393), .CLK (clk), .R (rst)) ;
    mux21_ni ix17394 (.Y (nx17393), .A0 (camera_module_cache_ram_139__6), .A1 (
             nx35572), .S0 (nx34332)) ;
    dffr camera_module_cache_reg_ram_155__6 (.Q (camera_module_cache_ram_155__6)
         , .QB (\$dummy [212]), .D (nx17383), .CLK (clk), .R (rst)) ;
    mux21_ni ix17384 (.Y (nx17383), .A0 (camera_module_cache_ram_155__6), .A1 (
             nx35572), .S0 (nx34328)) ;
    aoi22 ix24416 (.Y (nx24415), .A0 (camera_module_cache_ram_187__6), .A1 (
          nx36210), .B0 (camera_module_cache_ram_171__6), .B1 (nx36250)) ;
    dffr camera_module_cache_reg_ram_187__6 (.Q (camera_module_cache_ram_187__6)
         , .QB (\$dummy [213]), .D (nx17363), .CLK (clk), .R (rst)) ;
    mux21_ni ix17364 (.Y (nx17363), .A0 (camera_module_cache_ram_187__6), .A1 (
             nx35572), .S0 (nx34320)) ;
    dffr camera_module_cache_reg_ram_171__6 (.Q (camera_module_cache_ram_171__6)
         , .QB (\$dummy [214]), .D (nx17373), .CLK (clk), .R (rst)) ;
    mux21_ni ix17374 (.Y (nx17373), .A0 (camera_module_cache_ram_171__6), .A1 (
             nx35572), .S0 (nx34324)) ;
    aoi22 ix24429 (.Y (nx24428), .A0 (camera_module_cache_ram_203__6), .A1 (
          nx36290), .B0 (camera_module_cache_ram_219__6), .B1 (nx36330)) ;
    dffr camera_module_cache_reg_ram_203__6 (.Q (camera_module_cache_ram_203__6)
         , .QB (\$dummy [215]), .D (nx17353), .CLK (clk), .R (rst)) ;
    mux21_ni ix17354 (.Y (nx17353), .A0 (camera_module_cache_ram_203__6), .A1 (
             nx35572), .S0 (nx34316)) ;
    dffr camera_module_cache_reg_ram_219__6 (.Q (camera_module_cache_ram_219__6)
         , .QB (\$dummy [216]), .D (nx17343), .CLK (clk), .R (rst)) ;
    mux21_ni ix17344 (.Y (nx17343), .A0 (camera_module_cache_ram_219__6), .A1 (
             nx35574), .S0 (nx34312)) ;
    aoi22 ix24441 (.Y (nx24440), .A0 (camera_module_cache_ram_235__6), .A1 (
          nx36370), .B0 (camera_module_cache_ram_251__6), .B1 (nx36410)) ;
    dffr camera_module_cache_reg_ram_235__6 (.Q (camera_module_cache_ram_235__6)
         , .QB (\$dummy [217]), .D (nx17333), .CLK (clk), .R (rst)) ;
    mux21_ni ix17334 (.Y (nx17333), .A0 (camera_module_cache_ram_235__6), .A1 (
             nx35574), .S0 (nx34308)) ;
    dffr camera_module_cache_reg_ram_251__6 (.Q (camera_module_cache_ram_251__6)
         , .QB (\$dummy [218]), .D (nx17323), .CLK (clk), .R (rst)) ;
    mux21_ni ix17324 (.Y (nx17323), .A0 (camera_module_cache_ram_251__6), .A1 (
             nx35574), .S0 (nx34304)) ;
    nand04 ix20625 (.Y (nx20624), .A0 (nx24455), .A1 (nx24572), .A2 (nx24686), .A3 (
           nx24801)) ;
    oai21 ix24456 (.Y (nx24455), .A0 (nx20614), .A1 (nx20536), .B0 (nx36506)) ;
    nand04 ix20615 (.Y (nx20614), .A0 (nx24459), .A1 (nx24477), .A2 (nx24490), .A3 (
           nx24503)) ;
    aoi22 ix24460 (.Y (nx24459), .A0 (camera_module_cache_ram_12__6), .A1 (
          nx35810), .B0 (camera_module_cache_ram_28__6), .B1 (nx35850)) ;
    dffr camera_module_cache_reg_ram_12__6 (.Q (camera_module_cache_ram_12__6), 
         .QB (\$dummy [219]), .D (nx17313), .CLK (clk), .R (rst)) ;
    mux21_ni ix17314 (.Y (nx17313), .A0 (nx35574), .A1 (
             camera_module_cache_ram_12__6), .S0 (nx36496)) ;
    nand02 ix913 (.Y (nx912), .A0 (nx906), .A1 (nx880)) ;
    dffr camera_module_cache_reg_ram_28__6 (.Q (camera_module_cache_ram_28__6), 
         .QB (\$dummy [220]), .D (nx17303), .CLK (clk), .R (rst)) ;
    mux21_ni ix17304 (.Y (nx17303), .A0 (nx35574), .A1 (
             camera_module_cache_ram_28__6), .S0 (nx36510)) ;
    aoi22 ix24478 (.Y (nx24477), .A0 (camera_module_cache_ram_44__6), .A1 (
          nx35890), .B0 (camera_module_cache_ram_60__6), .B1 (nx35930)) ;
    dffr camera_module_cache_reg_ram_44__6 (.Q (camera_module_cache_ram_44__6), 
         .QB (\$dummy [221]), .D (nx17293), .CLK (clk), .R (rst)) ;
    mux21_ni ix17294 (.Y (nx17293), .A0 (nx35574), .A1 (
             camera_module_cache_ram_44__6), .S0 (nx36514)) ;
    dffr camera_module_cache_reg_ram_60__6 (.Q (camera_module_cache_ram_60__6), 
         .QB (\$dummy [222]), .D (nx17283), .CLK (clk), .R (rst)) ;
    mux21_ni ix17284 (.Y (nx17283), .A0 (nx35574), .A1 (
             camera_module_cache_ram_60__6), .S0 (nx36518)) ;
    aoi22 ix24491 (.Y (nx24490), .A0 (camera_module_cache_ram_76__6), .A1 (
          nx35970), .B0 (camera_module_cache_ram_92__6), .B1 (nx36010)) ;
    dffr camera_module_cache_reg_ram_76__6 (.Q (camera_module_cache_ram_76__6), 
         .QB (\$dummy [223]), .D (nx17273), .CLK (clk), .R (rst)) ;
    mux21_ni ix17274 (.Y (nx17273), .A0 (nx35576), .A1 (
             camera_module_cache_ram_76__6), .S0 (nx36522)) ;
    dffr camera_module_cache_reg_ram_92__6 (.Q (camera_module_cache_ram_92__6), 
         .QB (\$dummy [224]), .D (nx17263), .CLK (clk), .R (rst)) ;
    mux21_ni ix17264 (.Y (nx17263), .A0 (nx35576), .A1 (
             camera_module_cache_ram_92__6), .S0 (nx36526)) ;
    aoi22 ix24504 (.Y (nx24503), .A0 (camera_module_cache_ram_124__6), .A1 (
          nx36050), .B0 (camera_module_cache_ram_108__6), .B1 (nx36090)) ;
    dffr camera_module_cache_reg_ram_124__6 (.Q (camera_module_cache_ram_124__6)
         , .QB (\$dummy [225]), .D (nx17243), .CLK (clk), .R (rst)) ;
    mux21_ni ix17244 (.Y (nx17243), .A0 (nx35576), .A1 (
             camera_module_cache_ram_124__6), .S0 (nx36530)) ;
    dffr camera_module_cache_reg_ram_108__6 (.Q (camera_module_cache_ram_108__6)
         , .QB (\$dummy [226]), .D (nx17253), .CLK (clk), .R (rst)) ;
    mux21_ni ix17254 (.Y (nx17253), .A0 (nx35576), .A1 (
             camera_module_cache_ram_108__6), .S0 (nx36534)) ;
    nand04 ix20537 (.Y (nx20536), .A0 (nx24517), .A1 (nx24529), .A2 (nx24544), .A3 (
           nx24557)) ;
    aoi22 ix24518 (.Y (nx24517), .A0 (camera_module_cache_ram_140__6), .A1 (
          nx36130), .B0 (camera_module_cache_ram_156__6), .B1 (nx36170)) ;
    dffr camera_module_cache_reg_ram_140__6 (.Q (camera_module_cache_ram_140__6)
         , .QB (\$dummy [227]), .D (nx17233), .CLK (clk), .R (rst)) ;
    mux21_ni ix17234 (.Y (nx17233), .A0 (nx35576), .A1 (
             camera_module_cache_ram_140__6), .S0 (nx36538)) ;
    dffr camera_module_cache_reg_ram_156__6 (.Q (camera_module_cache_ram_156__6)
         , .QB (\$dummy [228]), .D (nx17223), .CLK (clk), .R (rst)) ;
    mux21_ni ix17224 (.Y (nx17223), .A0 (nx35576), .A1 (
             camera_module_cache_ram_156__6), .S0 (nx36542)) ;
    aoi22 ix24530 (.Y (nx24529), .A0 (camera_module_cache_ram_188__6), .A1 (
          nx36210), .B0 (camera_module_cache_ram_172__6), .B1 (nx36250)) ;
    dffr camera_module_cache_reg_ram_188__6 (.Q (camera_module_cache_ram_188__6)
         , .QB (\$dummy [229]), .D (nx17203), .CLK (clk), .R (rst)) ;
    mux21_ni ix17204 (.Y (nx17203), .A0 (nx35576), .A1 (
             camera_module_cache_ram_188__6), .S0 (nx36546)) ;
    dffr camera_module_cache_reg_ram_172__6 (.Q (camera_module_cache_ram_172__6)
         , .QB (\$dummy [230]), .D (nx17213), .CLK (clk), .R (rst)) ;
    mux21_ni ix17214 (.Y (nx17213), .A0 (nx35578), .A1 (
             camera_module_cache_ram_172__6), .S0 (nx36550)) ;
    aoi22 ix24545 (.Y (nx24544), .A0 (camera_module_cache_ram_204__6), .A1 (
          nx36290), .B0 (camera_module_cache_ram_220__6), .B1 (nx36330)) ;
    dffr camera_module_cache_reg_ram_204__6 (.Q (camera_module_cache_ram_204__6)
         , .QB (\$dummy [231]), .D (nx17193), .CLK (clk), .R (rst)) ;
    mux21_ni ix17194 (.Y (nx17193), .A0 (nx35578), .A1 (
             camera_module_cache_ram_204__6), .S0 (nx36554)) ;
    dffr camera_module_cache_reg_ram_220__6 (.Q (camera_module_cache_ram_220__6)
         , .QB (\$dummy [232]), .D (nx17183), .CLK (clk), .R (rst)) ;
    mux21_ni ix17184 (.Y (nx17183), .A0 (nx35578), .A1 (
             camera_module_cache_ram_220__6), .S0 (nx36558)) ;
    aoi22 ix24558 (.Y (nx24557), .A0 (camera_module_cache_ram_236__6), .A1 (
          nx36370), .B0 (camera_module_cache_ram_252__6), .B1 (nx36410)) ;
    dffr camera_module_cache_reg_ram_236__6 (.Q (camera_module_cache_ram_236__6)
         , .QB (\$dummy [233]), .D (nx17173), .CLK (clk), .R (rst)) ;
    mux21_ni ix17174 (.Y (nx17173), .A0 (nx35578), .A1 (
             camera_module_cache_ram_236__6), .S0 (nx36562)) ;
    dffr camera_module_cache_reg_ram_252__6 (.Q (camera_module_cache_ram_252__6)
         , .QB (\$dummy [234]), .D (nx17163), .CLK (clk), .R (rst)) ;
    mux21_ni ix17164 (.Y (nx17163), .A0 (nx35578), .A1 (
             camera_module_cache_ram_252__6), .S0 (nx36566)) ;
    oai21 ix24573 (.Y (nx24572), .A0 (nx20452), .A1 (nx20374), .B0 (nx36580)) ;
    nand04 ix20453 (.Y (nx20452), .A0 (nx24575), .A1 (nx24592), .A2 (nx24605), .A3 (
           nx24619)) ;
    aoi22 ix24576 (.Y (nx24575), .A0 (camera_module_cache_ram_13__6), .A1 (
          nx35812), .B0 (camera_module_cache_ram_29__6), .B1 (nx35852)) ;
    dffr camera_module_cache_reg_ram_13__6 (.Q (camera_module_cache_ram_13__6), 
         .QB (\$dummy [235]), .D (nx17153), .CLK (clk), .R (rst)) ;
    mux21_ni ix17154 (.Y (nx17153), .A0 (nx35578), .A1 (
             camera_module_cache_ram_13__6), .S0 (nx36570)) ;
    dffr camera_module_cache_reg_ram_29__6 (.Q (camera_module_cache_ram_29__6), 
         .QB (\$dummy [236]), .D (nx17143), .CLK (clk), .R (rst)) ;
    mux21_ni ix17144 (.Y (nx17143), .A0 (nx35578), .A1 (
             camera_module_cache_ram_29__6), .S0 (nx36584)) ;
    aoi22 ix24593 (.Y (nx24592), .A0 (camera_module_cache_ram_45__6), .A1 (
          nx35892), .B0 (camera_module_cache_ram_61__6), .B1 (nx35932)) ;
    dffr camera_module_cache_reg_ram_45__6 (.Q (camera_module_cache_ram_45__6), 
         .QB (\$dummy [237]), .D (nx17133), .CLK (clk), .R (rst)) ;
    mux21_ni ix17134 (.Y (nx17133), .A0 (nx35580), .A1 (
             camera_module_cache_ram_45__6), .S0 (nx36588)) ;
    dffr camera_module_cache_reg_ram_61__6 (.Q (camera_module_cache_ram_61__6), 
         .QB (\$dummy [238]), .D (nx17123), .CLK (clk), .R (rst)) ;
    mux21_ni ix17124 (.Y (nx17123), .A0 (nx35580), .A1 (
             camera_module_cache_ram_61__6), .S0 (nx36592)) ;
    aoi22 ix24606 (.Y (nx24605), .A0 (camera_module_cache_ram_77__6), .A1 (
          nx35972), .B0 (camera_module_cache_ram_93__6), .B1 (nx36012)) ;
    dffr camera_module_cache_reg_ram_77__6 (.Q (camera_module_cache_ram_77__6), 
         .QB (\$dummy [239]), .D (nx17113), .CLK (clk), .R (rst)) ;
    mux21_ni ix17114 (.Y (nx17113), .A0 (nx35580), .A1 (
             camera_module_cache_ram_77__6), .S0 (nx36596)) ;
    dffr camera_module_cache_reg_ram_93__6 (.Q (camera_module_cache_ram_93__6), 
         .QB (\$dummy [240]), .D (nx17103), .CLK (clk), .R (rst)) ;
    mux21_ni ix17104 (.Y (nx17103), .A0 (nx35580), .A1 (
             camera_module_cache_ram_93__6), .S0 (nx36600)) ;
    aoi22 ix24620 (.Y (nx24619), .A0 (camera_module_cache_ram_125__6), .A1 (
          nx36052), .B0 (camera_module_cache_ram_109__6), .B1 (nx36092)) ;
    dffr camera_module_cache_reg_ram_125__6 (.Q (camera_module_cache_ram_125__6)
         , .QB (\$dummy [241]), .D (nx17083), .CLK (clk), .R (rst)) ;
    mux21_ni ix17084 (.Y (nx17083), .A0 (nx35580), .A1 (
             camera_module_cache_ram_125__6), .S0 (nx36604)) ;
    dffr camera_module_cache_reg_ram_109__6 (.Q (camera_module_cache_ram_109__6)
         , .QB (\$dummy [242]), .D (nx17093), .CLK (clk), .R (rst)) ;
    mux21_ni ix17094 (.Y (nx17093), .A0 (nx35580), .A1 (
             camera_module_cache_ram_109__6), .S0 (nx36608)) ;
    nand04 ix20375 (.Y (nx20374), .A0 (nx24633), .A1 (nx24645), .A2 (nx24659), .A3 (
           nx24672)) ;
    aoi22 ix24634 (.Y (nx24633), .A0 (camera_module_cache_ram_141__6), .A1 (
          nx36132), .B0 (camera_module_cache_ram_157__6), .B1 (nx36172)) ;
    dffr camera_module_cache_reg_ram_141__6 (.Q (camera_module_cache_ram_141__6)
         , .QB (\$dummy [243]), .D (nx17073), .CLK (clk), .R (rst)) ;
    mux21_ni ix17074 (.Y (nx17073), .A0 (nx35580), .A1 (
             camera_module_cache_ram_141__6), .S0 (nx36612)) ;
    dffr camera_module_cache_reg_ram_157__6 (.Q (camera_module_cache_ram_157__6)
         , .QB (\$dummy [244]), .D (nx17063), .CLK (clk), .R (rst)) ;
    mux21_ni ix17064 (.Y (nx17063), .A0 (nx35582), .A1 (
             camera_module_cache_ram_157__6), .S0 (nx36616)) ;
    aoi22 ix24646 (.Y (nx24645), .A0 (camera_module_cache_ram_189__6), .A1 (
          nx36212), .B0 (camera_module_cache_ram_173__6), .B1 (nx36252)) ;
    dffr camera_module_cache_reg_ram_189__6 (.Q (camera_module_cache_ram_189__6)
         , .QB (\$dummy [245]), .D (nx17043), .CLK (clk), .R (rst)) ;
    mux21_ni ix17044 (.Y (nx17043), .A0 (nx35582), .A1 (
             camera_module_cache_ram_189__6), .S0 (nx36620)) ;
    dffr camera_module_cache_reg_ram_173__6 (.Q (camera_module_cache_ram_173__6)
         , .QB (\$dummy [246]), .D (nx17053), .CLK (clk), .R (rst)) ;
    mux21_ni ix17054 (.Y (nx17053), .A0 (nx35582), .A1 (
             camera_module_cache_ram_173__6), .S0 (nx36624)) ;
    aoi22 ix24660 (.Y (nx24659), .A0 (camera_module_cache_ram_205__6), .A1 (
          nx36292), .B0 (camera_module_cache_ram_221__6), .B1 (nx36332)) ;
    dffr camera_module_cache_reg_ram_205__6 (.Q (camera_module_cache_ram_205__6)
         , .QB (\$dummy [247]), .D (nx17033), .CLK (clk), .R (rst)) ;
    mux21_ni ix17034 (.Y (nx17033), .A0 (nx35582), .A1 (
             camera_module_cache_ram_205__6), .S0 (nx36628)) ;
    dffr camera_module_cache_reg_ram_221__6 (.Q (camera_module_cache_ram_221__6)
         , .QB (\$dummy [248]), .D (nx17023), .CLK (clk), .R (rst)) ;
    mux21_ni ix17024 (.Y (nx17023), .A0 (nx35582), .A1 (
             camera_module_cache_ram_221__6), .S0 (nx36632)) ;
    aoi22 ix24673 (.Y (nx24672), .A0 (camera_module_cache_ram_237__6), .A1 (
          nx36372), .B0 (camera_module_cache_ram_253__6), .B1 (nx36412)) ;
    dffr camera_module_cache_reg_ram_237__6 (.Q (camera_module_cache_ram_237__6)
         , .QB (\$dummy [249]), .D (nx17013), .CLK (clk), .R (rst)) ;
    mux21_ni ix17014 (.Y (nx17013), .A0 (nx35582), .A1 (
             camera_module_cache_ram_237__6), .S0 (nx36636)) ;
    dffr camera_module_cache_reg_ram_253__6 (.Q (camera_module_cache_ram_253__6)
         , .QB (\$dummy [250]), .D (nx17003), .CLK (clk), .R (rst)) ;
    mux21_ni ix17004 (.Y (nx17003), .A0 (nx35582), .A1 (
             camera_module_cache_ram_253__6), .S0 (nx36640)) ;
    oai21 ix24687 (.Y (nx24686), .A0 (nx20288), .A1 (nx20210), .B0 (nx36654)) ;
    nand04 ix20289 (.Y (nx20288), .A0 (nx24689), .A1 (nx24707), .A2 (nx24720), .A3 (
           nx24733)) ;
    aoi22 ix24690 (.Y (nx24689), .A0 (camera_module_cache_ram_14__6), .A1 (
          nx35812), .B0 (camera_module_cache_ram_30__6), .B1 (nx35852)) ;
    dffr camera_module_cache_reg_ram_14__6 (.Q (camera_module_cache_ram_14__6), 
         .QB (\$dummy [251]), .D (nx16993), .CLK (clk), .R (rst)) ;
    mux21_ni ix16994 (.Y (nx16993), .A0 (nx35584), .A1 (
             camera_module_cache_ram_14__6), .S0 (nx36644)) ;
    dffr camera_module_cache_reg_ram_30__6 (.Q (camera_module_cache_ram_30__6), 
         .QB (\$dummy [252]), .D (nx16983), .CLK (clk), .R (rst)) ;
    mux21_ni ix16984 (.Y (nx16983), .A0 (nx35584), .A1 (
             camera_module_cache_ram_30__6), .S0 (nx36658)) ;
    aoi22 ix24708 (.Y (nx24707), .A0 (camera_module_cache_ram_46__6), .A1 (
          nx35892), .B0 (camera_module_cache_ram_62__6), .B1 (nx35932)) ;
    dffr camera_module_cache_reg_ram_46__6 (.Q (camera_module_cache_ram_46__6), 
         .QB (\$dummy [253]), .D (nx16973), .CLK (clk), .R (rst)) ;
    mux21_ni ix16974 (.Y (nx16973), .A0 (nx35584), .A1 (
             camera_module_cache_ram_46__6), .S0 (nx36662)) ;
    dffr camera_module_cache_reg_ram_62__6 (.Q (camera_module_cache_ram_62__6), 
         .QB (\$dummy [254]), .D (nx16963), .CLK (clk), .R (rst)) ;
    mux21_ni ix16964 (.Y (nx16963), .A0 (nx35584), .A1 (
             camera_module_cache_ram_62__6), .S0 (nx36666)) ;
    aoi22 ix24721 (.Y (nx24720), .A0 (camera_module_cache_ram_78__6), .A1 (
          nx35972), .B0 (camera_module_cache_ram_94__6), .B1 (nx36012)) ;
    dffr camera_module_cache_reg_ram_78__6 (.Q (camera_module_cache_ram_78__6), 
         .QB (\$dummy [255]), .D (nx16953), .CLK (clk), .R (rst)) ;
    mux21_ni ix16954 (.Y (nx16953), .A0 (nx35584), .A1 (
             camera_module_cache_ram_78__6), .S0 (nx36670)) ;
    dffr camera_module_cache_reg_ram_94__6 (.Q (camera_module_cache_ram_94__6), 
         .QB (\$dummy [256]), .D (nx16943), .CLK (clk), .R (rst)) ;
    mux21_ni ix16944 (.Y (nx16943), .A0 (nx35584), .A1 (
             camera_module_cache_ram_94__6), .S0 (nx36674)) ;
    aoi22 ix24734 (.Y (nx24733), .A0 (camera_module_cache_ram_126__6), .A1 (
          nx36052), .B0 (camera_module_cache_ram_110__6), .B1 (nx36092)) ;
    dffr camera_module_cache_reg_ram_126__6 (.Q (camera_module_cache_ram_126__6)
         , .QB (\$dummy [257]), .D (nx16923), .CLK (clk), .R (rst)) ;
    mux21_ni ix16924 (.Y (nx16923), .A0 (nx35584), .A1 (
             camera_module_cache_ram_126__6), .S0 (nx36678)) ;
    dffr camera_module_cache_reg_ram_110__6 (.Q (camera_module_cache_ram_110__6)
         , .QB (\$dummy [258]), .D (nx16933), .CLK (clk), .R (rst)) ;
    mux21_ni ix16934 (.Y (nx16933), .A0 (nx35586), .A1 (
             camera_module_cache_ram_110__6), .S0 (nx36682)) ;
    nand04 ix20211 (.Y (nx20210), .A0 (nx24747), .A1 (nx24760), .A2 (nx24774), .A3 (
           nx24788)) ;
    aoi22 ix24748 (.Y (nx24747), .A0 (camera_module_cache_ram_142__6), .A1 (
          nx36132), .B0 (camera_module_cache_ram_158__6), .B1 (nx36172)) ;
    dffr camera_module_cache_reg_ram_142__6 (.Q (camera_module_cache_ram_142__6)
         , .QB (\$dummy [259]), .D (nx16913), .CLK (clk), .R (rst)) ;
    mux21_ni ix16914 (.Y (nx16913), .A0 (nx35586), .A1 (
             camera_module_cache_ram_142__6), .S0 (nx36686)) ;
    dffr camera_module_cache_reg_ram_158__6 (.Q (camera_module_cache_ram_158__6)
         , .QB (\$dummy [260]), .D (nx16903), .CLK (clk), .R (rst)) ;
    mux21_ni ix16904 (.Y (nx16903), .A0 (nx35586), .A1 (
             camera_module_cache_ram_158__6), .S0 (nx36690)) ;
    aoi22 ix24761 (.Y (nx24760), .A0 (camera_module_cache_ram_190__6), .A1 (
          nx36212), .B0 (camera_module_cache_ram_174__6), .B1 (nx36252)) ;
    dffr camera_module_cache_reg_ram_190__6 (.Q (camera_module_cache_ram_190__6)
         , .QB (\$dummy [261]), .D (nx16883), .CLK (clk), .R (rst)) ;
    mux21_ni ix16884 (.Y (nx16883), .A0 (nx35586), .A1 (
             camera_module_cache_ram_190__6), .S0 (nx36694)) ;
    dffr camera_module_cache_reg_ram_174__6 (.Q (camera_module_cache_ram_174__6)
         , .QB (\$dummy [262]), .D (nx16893), .CLK (clk), .R (rst)) ;
    mux21_ni ix16894 (.Y (nx16893), .A0 (nx35586), .A1 (
             camera_module_cache_ram_174__6), .S0 (nx36698)) ;
    aoi22 ix24775 (.Y (nx24774), .A0 (camera_module_cache_ram_206__6), .A1 (
          nx36292), .B0 (camera_module_cache_ram_222__6), .B1 (nx36332)) ;
    dffr camera_module_cache_reg_ram_206__6 (.Q (camera_module_cache_ram_206__6)
         , .QB (\$dummy [263]), .D (nx16873), .CLK (clk), .R (rst)) ;
    mux21_ni ix16874 (.Y (nx16873), .A0 (nx35586), .A1 (
             camera_module_cache_ram_206__6), .S0 (nx36702)) ;
    dffr camera_module_cache_reg_ram_222__6 (.Q (camera_module_cache_ram_222__6)
         , .QB (\$dummy [264]), .D (nx16863), .CLK (clk), .R (rst)) ;
    mux21_ni ix16864 (.Y (nx16863), .A0 (nx35586), .A1 (
             camera_module_cache_ram_222__6), .S0 (nx36706)) ;
    aoi22 ix24789 (.Y (nx24788), .A0 (camera_module_cache_ram_238__6), .A1 (
          nx36372), .B0 (camera_module_cache_ram_254__6), .B1 (nx36412)) ;
    dffr camera_module_cache_reg_ram_238__6 (.Q (camera_module_cache_ram_238__6)
         , .QB (\$dummy [265]), .D (nx16853), .CLK (clk), .R (rst)) ;
    mux21_ni ix16854 (.Y (nx16853), .A0 (nx35588), .A1 (
             camera_module_cache_ram_238__6), .S0 (nx36710)) ;
    dffr camera_module_cache_reg_ram_254__6 (.Q (camera_module_cache_ram_254__6)
         , .QB (\$dummy [266]), .D (nx16843), .CLK (clk), .R (rst)) ;
    mux21_ni ix16844 (.Y (nx16843), .A0 (nx35588), .A1 (
             camera_module_cache_ram_254__6), .S0 (nx36714)) ;
    oai21 ix24802 (.Y (nx24801), .A0 (nx20126), .A1 (nx20048), .B0 (nx36728)) ;
    nand04 ix20127 (.Y (nx20126), .A0 (nx24805), .A1 (nx24819), .A2 (nx24834), .A3 (
           nx24848)) ;
    aoi22 ix24806 (.Y (nx24805), .A0 (camera_module_cache_ram_15__6), .A1 (
          nx35812), .B0 (camera_module_cache_ram_31__6), .B1 (nx35852)) ;
    dffr camera_module_cache_reg_ram_15__6 (.Q (camera_module_cache_ram_15__6), 
         .QB (\$dummy [267]), .D (nx16833), .CLK (clk), .R (rst)) ;
    mux21_ni ix16834 (.Y (nx16833), .A0 (nx35588), .A1 (
             camera_module_cache_ram_15__6), .S0 (nx36718)) ;
    nor02_2x ix24812 (.Y (nx24811), .A0 (nx912), .A1 (nx842)) ;
    dffr camera_module_cache_reg_ram_31__6 (.Q (camera_module_cache_ram_31__6), 
         .QB (\$dummy [268]), .D (nx16823), .CLK (clk), .R (rst)) ;
    mux21_ni ix16824 (.Y (nx16823), .A0 (nx35588), .A1 (
             camera_module_cache_ram_31__6), .S0 (nx36732)) ;
    aoi22 ix24820 (.Y (nx24819), .A0 (camera_module_cache_ram_47__6), .A1 (
          nx35892), .B0 (camera_module_cache_ram_63__6), .B1 (nx35932)) ;
    dffr camera_module_cache_reg_ram_47__6 (.Q (camera_module_cache_ram_47__6), 
         .QB (\$dummy [269]), .D (nx16813), .CLK (clk), .R (rst)) ;
    mux21_ni ix16814 (.Y (nx16813), .A0 (nx35588), .A1 (
             camera_module_cache_ram_47__6), .S0 (nx36736)) ;
    dffr camera_module_cache_reg_ram_63__6 (.Q (camera_module_cache_ram_63__6), 
         .QB (\$dummy [270]), .D (nx16803), .CLK (clk), .R (rst)) ;
    mux21_ni ix16804 (.Y (nx16803), .A0 (nx35588), .A1 (
             camera_module_cache_ram_63__6), .S0 (nx36740)) ;
    aoi22 ix24835 (.Y (nx24834), .A0 (camera_module_cache_ram_79__6), .A1 (
          nx35972), .B0 (camera_module_cache_ram_95__6), .B1 (nx36012)) ;
    dffr camera_module_cache_reg_ram_79__6 (.Q (camera_module_cache_ram_79__6), 
         .QB (\$dummy [271]), .D (nx16793), .CLK (clk), .R (rst)) ;
    mux21_ni ix16794 (.Y (nx16793), .A0 (nx35588), .A1 (
             camera_module_cache_ram_79__6), .S0 (nx36744)) ;
    dffr camera_module_cache_reg_ram_95__6 (.Q (camera_module_cache_ram_95__6), 
         .QB (\$dummy [272]), .D (nx16783), .CLK (clk), .R (rst)) ;
    mux21_ni ix16784 (.Y (nx16783), .A0 (nx35590), .A1 (
             camera_module_cache_ram_95__6), .S0 (nx36748)) ;
    aoi22 ix24849 (.Y (nx24848), .A0 (camera_module_cache_ram_127__6), .A1 (
          nx36052), .B0 (camera_module_cache_ram_111__6), .B1 (nx36092)) ;
    dffr camera_module_cache_reg_ram_127__6 (.Q (camera_module_cache_ram_127__6)
         , .QB (\$dummy [273]), .D (nx16763), .CLK (clk), .R (rst)) ;
    mux21_ni ix16764 (.Y (nx16763), .A0 (nx35590), .A1 (
             camera_module_cache_ram_127__6), .S0 (nx36752)) ;
    dffr camera_module_cache_reg_ram_111__6 (.Q (camera_module_cache_ram_111__6)
         , .QB (\$dummy [274]), .D (nx16773), .CLK (clk), .R (rst)) ;
    mux21_ni ix16774 (.Y (nx16773), .A0 (nx35590), .A1 (
             camera_module_cache_ram_111__6), .S0 (nx36756)) ;
    nand04 ix20049 (.Y (nx20048), .A0 (nx24863), .A1 (nx24877), .A2 (nx24890), .A3 (
           nx24903)) ;
    aoi22 ix24864 (.Y (nx24863), .A0 (camera_module_cache_ram_143__6), .A1 (
          nx36132), .B0 (camera_module_cache_ram_159__6), .B1 (nx36172)) ;
    dffr camera_module_cache_reg_ram_143__6 (.Q (camera_module_cache_ram_143__6)
         , .QB (\$dummy [275]), .D (nx16753), .CLK (clk), .R (rst)) ;
    mux21_ni ix16754 (.Y (nx16753), .A0 (nx35590), .A1 (
             camera_module_cache_ram_143__6), .S0 (nx36760)) ;
    dffr camera_module_cache_reg_ram_159__6 (.Q (camera_module_cache_ram_159__6)
         , .QB (\$dummy [276]), .D (nx16743), .CLK (clk), .R (rst)) ;
    mux21_ni ix16744 (.Y (nx16743), .A0 (nx35590), .A1 (
             camera_module_cache_ram_159__6), .S0 (nx36764)) ;
    aoi22 ix24878 (.Y (nx24877), .A0 (camera_module_cache_ram_191__6), .A1 (
          nx36212), .B0 (camera_module_cache_ram_175__6), .B1 (nx36252)) ;
    dffr camera_module_cache_reg_ram_191__6 (.Q (camera_module_cache_ram_191__6)
         , .QB (\$dummy [277]), .D (nx16723), .CLK (clk), .R (rst)) ;
    mux21_ni ix16724 (.Y (nx16723), .A0 (nx35590), .A1 (
             camera_module_cache_ram_191__6), .S0 (nx36768)) ;
    dffr camera_module_cache_reg_ram_175__6 (.Q (camera_module_cache_ram_175__6)
         , .QB (\$dummy [278]), .D (nx16733), .CLK (clk), .R (rst)) ;
    mux21_ni ix16734 (.Y (nx16733), .A0 (nx35590), .A1 (
             camera_module_cache_ram_175__6), .S0 (nx36772)) ;
    aoi22 ix24891 (.Y (nx24890), .A0 (camera_module_cache_ram_207__6), .A1 (
          nx36292), .B0 (camera_module_cache_ram_223__6), .B1 (nx36332)) ;
    dffr camera_module_cache_reg_ram_207__6 (.Q (camera_module_cache_ram_207__6)
         , .QB (\$dummy [279]), .D (nx16713), .CLK (clk), .R (rst)) ;
    mux21_ni ix16714 (.Y (nx16713), .A0 (nx35592), .A1 (
             camera_module_cache_ram_207__6), .S0 (nx36776)) ;
    dffr camera_module_cache_reg_ram_223__6 (.Q (camera_module_cache_ram_223__6)
         , .QB (\$dummy [280]), .D (nx16703), .CLK (clk), .R (rst)) ;
    mux21_ni ix16704 (.Y (nx16703), .A0 (nx35592), .A1 (
             camera_module_cache_ram_223__6), .S0 (nx36780)) ;
    aoi22 ix24904 (.Y (nx24903), .A0 (camera_module_cache_ram_239__6), .A1 (
          nx36372), .B0 (camera_module_cache_ram_255__6), .B1 (nx36412)) ;
    dffr camera_module_cache_reg_ram_239__6 (.Q (camera_module_cache_ram_239__6)
         , .QB (\$dummy [281]), .D (nx16693), .CLK (clk), .R (rst)) ;
    mux21_ni ix16694 (.Y (nx16693), .A0 (nx35592), .A1 (
             camera_module_cache_ram_239__6), .S0 (nx36784)) ;
    dffr camera_module_cache_reg_ram_255__6 (.Q (camera_module_cache_ram_255__6)
         , .QB (\$dummy [282]), .D (nx16683), .CLK (clk), .R (rst)) ;
    mux21_ni ix16684 (.Y (nx16683), .A0 (nx35592), .A1 (
             camera_module_cache_ram_255__6), .S0 (nx36788)) ;
    aoi21 ix24919 (.Y (nx24918), .A0 (nx35806), .A1 (nx770), .B0 (nx738)) ;
    nand03 ix771 (.Y (nx770), .A0 (nx24921), .A1 (nx37082), .A2 (nx24925)) ;
    aoi21 ix24926 (.Y (nx24925), .A0 (camera_module_algo_module_address_value_3)
          , .A1 (nx23021), .B0 (nx752)) ;
    aoi21 ix740 (.Y (nx738), .A0 (nx24930), .A1 (nx24933), .B0 (nx35806)) ;
    aoi21 ix24931 (.Y (nx24930), .A0 (nx37094), .A1 (nx622), .B0 (nx37082)) ;
    nor04 ix623 (.Y (nx622), .A0 (camera_module_algo_module_address_value_7), .A1 (
          camera_module_algo_module_address_value_6), .A2 (
          camera_module_algo_module_address_value_5), .A3 (
          camera_module_algo_module_address_value_4)) ;
    mux21_ni ix24934 (.Y (nx24933), .A0 (nx37094), .A1 (nx622), .S0 (nx24935)) ;
    nand04 ix24936 (.Y (nx24935), .A0 (camera_module_algo_module_address_value_7
           ), .A1 (camera_module_algo_module_address_value_6), .A2 (
           camera_module_algo_module_address_value_5), .A3 (
           camera_module_algo_module_address_value_4)) ;
    oai22 ix19851 (.Y (nx19850), .A0 (nx24939), .A1 (nx31101), .B0 (nx32240), .B1 (
          nx19826)) ;
    aoi22 ix24940 (.Y (nx24939), .A0 (camera_module_algo_module_pixel_value_4), 
          .A1 (nx24945), .B0 (nx14302), .B1 (nx17068)) ;
    dff camera_module_algo_module_pixel_reg_reg_q_4 (.Q (
        camera_module_algo_module_pixel_value_4), .QB (\$dummy [283]), .D (
        nx14103), .CLK (clk)) ;
    mux21_ni ix14104 (.Y (nx14103), .A0 (nx17060), .A1 (
             camera_module_algo_module_pixel_value_4), .S0 (nx37152)) ;
    mux21_ni ix24946 (.Y (nx24945), .A0 (nx24947), .A1 (nx35674), .S0 (nx36792)
             ) ;
    nor04 ix24948 (.Y (nx24947), .A0 (nx17040), .A1 (nx16386), .A2 (nx15730), .A3 (
          nx15076)) ;
    nand04 ix17041 (.Y (nx17040), .A0 (nx24951), .A1 (nx25074), .A2 (nx25149), .A3 (
           nx25227)) ;
    oai21 ix24952 (.Y (nx24951), .A0 (nx17030), .A1 (nx16952), .B0 (nx36448)) ;
    nand04 ix17031 (.Y (nx17030), .A0 (nx24954), .A1 (nx25009), .A2 (nx25017), .A3 (
           nx25027)) ;
    aoi22 ix24955 (.Y (nx24954), .A0 (camera_module_cache_ram_0__4), .A1 (
          nx35812), .B0 (camera_module_cache_ram_16__4), .B1 (nx35852)) ;
    dffr camera_module_cache_reg_ram_0__4 (.Q (camera_module_cache_ram_0__4), .QB (
         \$dummy [284]), .D (nx14093), .CLK (clk), .R (rst)) ;
    mux21_ni ix14094 (.Y (nx14093), .A0 (camera_module_cache_ram_0__4), .A1 (
             nx35368), .S0 (nx35134)) ;
    oai221 ix14423 (.Y (nx14422), .A0 (nx34072), .A1 (nx24960), .B0 (nx24979), .B1 (
           nx35712), .C0 (nx24983)) ;
    tri01 nvm_module_tri_dataout_124 (.Y (nvm_data_124), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_116 (.Y (nvm_data_116), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_108 (.Y (nvm_data_108), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_100 (.Y (nvm_data_100), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_92 (.Y (nvm_data_92), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_84 (.Y (nvm_data_84), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_76 (.Y (nvm_data_76), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_68 (.Y (nvm_data_68), .A (nx22549), .E (
          nvm_module_GND0)) ;
    inv01 ix24980 (.Y (nx24979), .A (nvm_data_4)) ;
    tri01 nvm_module_tri_dataout_4 (.Y (nvm_data_4), .A (nx22549), .E (
          nvm_module_GND0)) ;
    nand02 ix24984 (.Y (nx24983), .A0 (nx34074), .A1 (nx14356)) ;
    tri01 nvm_module_tri_dataout_60 (.Y (nvm_data_60), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_52 (.Y (nvm_data_52), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_44 (.Y (nvm_data_44), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_36 (.Y (nvm_data_36), .A (nx22549), .E (
          nvm_module_GND0)) ;
    oai22 ix14325 (.Y (nx14324), .A0 (nx34100), .A1 (nx24997), .B0 (nx34082), .B1 (
          nx25001)) ;
    tri01 nvm_module_tri_dataout_28 (.Y (nvm_data_28), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_20 (.Y (nvm_data_20), .A (nx22549), .E (
          nvm_module_GND0)) ;
    nand02 ix25002 (.Y (nx25001), .A0 (nvm_data_12), .A1 (nx34100)) ;
    tri01 nvm_module_tri_dataout_12 (.Y (nvm_data_12), .A (nx22549), .E (
          nvm_module_GND0)) ;
    dffr camera_module_cache_reg_ram_16__4 (.Q (camera_module_cache_ram_16__4), 
         .QB (\$dummy [285]), .D (nx14083), .CLK (clk), .R (rst)) ;
    mux21_ni ix14084 (.Y (nx14083), .A0 (camera_module_cache_ram_16__4), .A1 (
             nx35368), .S0 (nx35130)) ;
    aoi22 ix25010 (.Y (nx25009), .A0 (camera_module_cache_ram_32__4), .A1 (
          nx35892), .B0 (camera_module_cache_ram_48__4), .B1 (nx35932)) ;
    dffr camera_module_cache_reg_ram_32__4 (.Q (camera_module_cache_ram_32__4), 
         .QB (\$dummy [286]), .D (nx14073), .CLK (clk), .R (rst)) ;
    mux21_ni ix14074 (.Y (nx14073), .A0 (camera_module_cache_ram_32__4), .A1 (
             nx35368), .S0 (nx35126)) ;
    dffr camera_module_cache_reg_ram_48__4 (.Q (camera_module_cache_ram_48__4), 
         .QB (\$dummy [287]), .D (nx14063), .CLK (clk), .R (rst)) ;
    mux21_ni ix14064 (.Y (nx14063), .A0 (camera_module_cache_ram_48__4), .A1 (
             nx35368), .S0 (nx35122)) ;
    aoi22 ix25018 (.Y (nx25017), .A0 (camera_module_cache_ram_64__4), .A1 (
          nx35972), .B0 (camera_module_cache_ram_80__4), .B1 (nx36012)) ;
    dffr camera_module_cache_reg_ram_64__4 (.Q (camera_module_cache_ram_64__4), 
         .QB (\$dummy [288]), .D (nx14053), .CLK (clk), .R (rst)) ;
    mux21_ni ix14054 (.Y (nx14053), .A0 (camera_module_cache_ram_64__4), .A1 (
             nx35368), .S0 (nx35118)) ;
    dffr camera_module_cache_reg_ram_80__4 (.Q (camera_module_cache_ram_80__4), 
         .QB (\$dummy [289]), .D (nx14043), .CLK (clk), .R (rst)) ;
    mux21_ni ix14044 (.Y (nx14043), .A0 (camera_module_cache_ram_80__4), .A1 (
             nx35368), .S0 (nx35114)) ;
    aoi22 ix25028 (.Y (nx25027), .A0 (camera_module_cache_ram_112__4), .A1 (
          nx36052), .B0 (camera_module_cache_ram_96__4), .B1 (nx36092)) ;
    dffr camera_module_cache_reg_ram_112__4 (.Q (camera_module_cache_ram_112__4)
         , .QB (\$dummy [290]), .D (nx14023), .CLK (clk), .R (rst)) ;
    mux21_ni ix14024 (.Y (nx14023), .A0 (camera_module_cache_ram_112__4), .A1 (
             nx35368), .S0 (nx35106)) ;
    dffr camera_module_cache_reg_ram_96__4 (.Q (camera_module_cache_ram_96__4), 
         .QB (\$dummy [291]), .D (nx14033), .CLK (clk), .R (rst)) ;
    mux21_ni ix14034 (.Y (nx14033), .A0 (camera_module_cache_ram_96__4), .A1 (
             nx35370), .S0 (nx35110)) ;
    nand04 ix16953 (.Y (nx16952), .A0 (nx25039), .A1 (nx25047), .A2 (nx25056), .A3 (
           nx25065)) ;
    aoi22 ix25040 (.Y (nx25039), .A0 (camera_module_cache_ram_128__4), .A1 (
          nx36132), .B0 (camera_module_cache_ram_144__4), .B1 (nx36172)) ;
    dffr camera_module_cache_reg_ram_128__4 (.Q (camera_module_cache_ram_128__4)
         , .QB (\$dummy [292]), .D (nx14013), .CLK (clk), .R (rst)) ;
    mux21_ni ix14014 (.Y (nx14013), .A0 (camera_module_cache_ram_128__4), .A1 (
             nx35370), .S0 (nx35102)) ;
    dffr camera_module_cache_reg_ram_144__4 (.Q (camera_module_cache_ram_144__4)
         , .QB (\$dummy [293]), .D (nx14003), .CLK (clk), .R (rst)) ;
    mux21_ni ix14004 (.Y (nx14003), .A0 (camera_module_cache_ram_144__4), .A1 (
             nx35370), .S0 (nx35098)) ;
    aoi22 ix25048 (.Y (nx25047), .A0 (camera_module_cache_ram_176__4), .A1 (
          nx36212), .B0 (camera_module_cache_ram_160__4), .B1 (nx36252)) ;
    dffr camera_module_cache_reg_ram_176__4 (.Q (camera_module_cache_ram_176__4)
         , .QB (\$dummy [294]), .D (nx13983), .CLK (clk), .R (rst)) ;
    mux21_ni ix13984 (.Y (nx13983), .A0 (camera_module_cache_ram_176__4), .A1 (
             nx35370), .S0 (nx35090)) ;
    dffr camera_module_cache_reg_ram_160__4 (.Q (camera_module_cache_ram_160__4)
         , .QB (\$dummy [295]), .D (nx13993), .CLK (clk), .R (rst)) ;
    mux21_ni ix13994 (.Y (nx13993), .A0 (camera_module_cache_ram_160__4), .A1 (
             nx35370), .S0 (nx35094)) ;
    aoi22 ix25057 (.Y (nx25056), .A0 (camera_module_cache_ram_192__4), .A1 (
          nx36292), .B0 (camera_module_cache_ram_208__4), .B1 (nx36332)) ;
    dffr camera_module_cache_reg_ram_192__4 (.Q (camera_module_cache_ram_192__4)
         , .QB (\$dummy [296]), .D (nx13973), .CLK (clk), .R (rst)) ;
    mux21_ni ix13974 (.Y (nx13973), .A0 (camera_module_cache_ram_192__4), .A1 (
             nx35370), .S0 (nx35086)) ;
    dffr camera_module_cache_reg_ram_208__4 (.Q (camera_module_cache_ram_208__4)
         , .QB (\$dummy [297]), .D (nx13963), .CLK (clk), .R (rst)) ;
    mux21_ni ix13964 (.Y (nx13963), .A0 (camera_module_cache_ram_208__4), .A1 (
             nx35370), .S0 (nx35082)) ;
    aoi22 ix25066 (.Y (nx25065), .A0 (camera_module_cache_ram_224__4), .A1 (
          nx36372), .B0 (camera_module_cache_ram_240__4), .B1 (nx36412)) ;
    dffr camera_module_cache_reg_ram_224__4 (.Q (camera_module_cache_ram_224__4)
         , .QB (\$dummy [298]), .D (nx13953), .CLK (clk), .R (rst)) ;
    mux21_ni ix13954 (.Y (nx13953), .A0 (camera_module_cache_ram_224__4), .A1 (
             nx35372), .S0 (nx35078)) ;
    dffr camera_module_cache_reg_ram_240__4 (.Q (camera_module_cache_ram_240__4)
         , .QB (\$dummy [299]), .D (nx13943), .CLK (clk), .R (rst)) ;
    mux21_ni ix13944 (.Y (nx13943), .A0 (camera_module_cache_ram_240__4), .A1 (
             nx35372), .S0 (nx35074)) ;
    oai21 ix25075 (.Y (nx25074), .A0 (nx16868), .A1 (nx16790), .B0 (nx36452)) ;
    nand04 ix16869 (.Y (nx16868), .A0 (nx25077), .A1 (nx25085), .A2 (nx25094), .A3 (
           nx25103)) ;
    aoi22 ix25078 (.Y (nx25077), .A0 (camera_module_cache_ram_1__4), .A1 (
          nx35814), .B0 (camera_module_cache_ram_17__4), .B1 (nx35854)) ;
    dffr camera_module_cache_reg_ram_1__4 (.Q (camera_module_cache_ram_1__4), .QB (
         \$dummy [300]), .D (nx13933), .CLK (clk), .R (rst)) ;
    mux21_ni ix13934 (.Y (nx13933), .A0 (camera_module_cache_ram_1__4), .A1 (
             nx35372), .S0 (nx35064)) ;
    dffr camera_module_cache_reg_ram_17__4 (.Q (camera_module_cache_ram_17__4), 
         .QB (\$dummy [301]), .D (nx13923), .CLK (clk), .R (rst)) ;
    mux21_ni ix13924 (.Y (nx13923), .A0 (camera_module_cache_ram_17__4), .A1 (
             nx35372), .S0 (nx35060)) ;
    aoi22 ix25086 (.Y (nx25085), .A0 (camera_module_cache_ram_33__4), .A1 (
          nx35894), .B0 (camera_module_cache_ram_49__4), .B1 (nx35934)) ;
    dffr camera_module_cache_reg_ram_33__4 (.Q (camera_module_cache_ram_33__4), 
         .QB (\$dummy [302]), .D (nx13913), .CLK (clk), .R (rst)) ;
    mux21_ni ix13914 (.Y (nx13913), .A0 (camera_module_cache_ram_33__4), .A1 (
             nx35372), .S0 (nx35056)) ;
    dffr camera_module_cache_reg_ram_49__4 (.Q (camera_module_cache_ram_49__4), 
         .QB (\$dummy [303]), .D (nx13903), .CLK (clk), .R (rst)) ;
    mux21_ni ix13904 (.Y (nx13903), .A0 (camera_module_cache_ram_49__4), .A1 (
             nx35372), .S0 (nx35052)) ;
    aoi22 ix25095 (.Y (nx25094), .A0 (camera_module_cache_ram_65__4), .A1 (
          nx35974), .B0 (camera_module_cache_ram_81__4), .B1 (nx36014)) ;
    dffr camera_module_cache_reg_ram_65__4 (.Q (camera_module_cache_ram_65__4), 
         .QB (\$dummy [304]), .D (nx13893), .CLK (clk), .R (rst)) ;
    mux21_ni ix13894 (.Y (nx13893), .A0 (camera_module_cache_ram_65__4), .A1 (
             nx35372), .S0 (nx35048)) ;
    dffr camera_module_cache_reg_ram_81__4 (.Q (camera_module_cache_ram_81__4), 
         .QB (\$dummy [305]), .D (nx13883), .CLK (clk), .R (rst)) ;
    mux21_ni ix13884 (.Y (nx13883), .A0 (camera_module_cache_ram_81__4), .A1 (
             nx35374), .S0 (nx35044)) ;
    aoi22 ix25104 (.Y (nx25103), .A0 (camera_module_cache_ram_113__4), .A1 (
          nx36054), .B0 (camera_module_cache_ram_97__4), .B1 (nx36094)) ;
    dffr camera_module_cache_reg_ram_113__4 (.Q (camera_module_cache_ram_113__4)
         , .QB (\$dummy [306]), .D (nx13863), .CLK (clk), .R (rst)) ;
    mux21_ni ix13864 (.Y (nx13863), .A0 (camera_module_cache_ram_113__4), .A1 (
             nx35374), .S0 (nx35036)) ;
    dffr camera_module_cache_reg_ram_97__4 (.Q (camera_module_cache_ram_97__4), 
         .QB (\$dummy [307]), .D (nx13873), .CLK (clk), .R (rst)) ;
    mux21_ni ix13874 (.Y (nx13873), .A0 (camera_module_cache_ram_97__4), .A1 (
             nx35374), .S0 (nx35040)) ;
    nand04 ix16791 (.Y (nx16790), .A0 (nx25113), .A1 (nx25122), .A2 (nx25131), .A3 (
           nx25140)) ;
    aoi22 ix25114 (.Y (nx25113), .A0 (camera_module_cache_ram_129__4), .A1 (
          nx36134), .B0 (camera_module_cache_ram_145__4), .B1 (nx36174)) ;
    dffr camera_module_cache_reg_ram_129__4 (.Q (camera_module_cache_ram_129__4)
         , .QB (\$dummy [308]), .D (nx13853), .CLK (clk), .R (rst)) ;
    mux21_ni ix13854 (.Y (nx13853), .A0 (camera_module_cache_ram_129__4), .A1 (
             nx35374), .S0 (nx35032)) ;
    dffr camera_module_cache_reg_ram_145__4 (.Q (camera_module_cache_ram_145__4)
         , .QB (\$dummy [309]), .D (nx13843), .CLK (clk), .R (rst)) ;
    mux21_ni ix13844 (.Y (nx13843), .A0 (camera_module_cache_ram_145__4), .A1 (
             nx35374), .S0 (nx35028)) ;
    aoi22 ix25123 (.Y (nx25122), .A0 (camera_module_cache_ram_177__4), .A1 (
          nx36214), .B0 (camera_module_cache_ram_161__4), .B1 (nx36254)) ;
    dffr camera_module_cache_reg_ram_177__4 (.Q (camera_module_cache_ram_177__4)
         , .QB (\$dummy [310]), .D (nx13823), .CLK (clk), .R (rst)) ;
    mux21_ni ix13824 (.Y (nx13823), .A0 (camera_module_cache_ram_177__4), .A1 (
             nx35374), .S0 (nx35020)) ;
    dffr camera_module_cache_reg_ram_161__4 (.Q (camera_module_cache_ram_161__4)
         , .QB (\$dummy [311]), .D (nx13833), .CLK (clk), .R (rst)) ;
    mux21_ni ix13834 (.Y (nx13833), .A0 (camera_module_cache_ram_161__4), .A1 (
             nx35374), .S0 (nx35024)) ;
    aoi22 ix25132 (.Y (nx25131), .A0 (camera_module_cache_ram_193__4), .A1 (
          nx36294), .B0 (camera_module_cache_ram_209__4), .B1 (nx36334)) ;
    dffr camera_module_cache_reg_ram_193__4 (.Q (camera_module_cache_ram_193__4)
         , .QB (\$dummy [312]), .D (nx13813), .CLK (clk), .R (rst)) ;
    mux21_ni ix13814 (.Y (nx13813), .A0 (camera_module_cache_ram_193__4), .A1 (
             nx35376), .S0 (nx35016)) ;
    dffr camera_module_cache_reg_ram_209__4 (.Q (camera_module_cache_ram_209__4)
         , .QB (\$dummy [313]), .D (nx13803), .CLK (clk), .R (rst)) ;
    mux21_ni ix13804 (.Y (nx13803), .A0 (camera_module_cache_ram_209__4), .A1 (
             nx35376), .S0 (nx35012)) ;
    aoi22 ix25141 (.Y (nx25140), .A0 (camera_module_cache_ram_225__4), .A1 (
          nx36374), .B0 (camera_module_cache_ram_241__4), .B1 (nx36414)) ;
    dffr camera_module_cache_reg_ram_225__4 (.Q (camera_module_cache_ram_225__4)
         , .QB (\$dummy [314]), .D (nx13793), .CLK (clk), .R (rst)) ;
    mux21_ni ix13794 (.Y (nx13793), .A0 (camera_module_cache_ram_225__4), .A1 (
             nx35376), .S0 (nx35008)) ;
    dffr camera_module_cache_reg_ram_241__4 (.Q (camera_module_cache_ram_241__4)
         , .QB (\$dummy [315]), .D (nx13783), .CLK (clk), .R (rst)) ;
    mux21_ni ix13784 (.Y (nx13783), .A0 (camera_module_cache_ram_241__4), .A1 (
             nx35376), .S0 (nx35004)) ;
    oai21 ix25150 (.Y (nx25149), .A0 (nx16704), .A1 (nx16626), .B0 (nx36456)) ;
    nand04 ix16705 (.Y (nx16704), .A0 (nx25153), .A1 (nx25162), .A2 (nx25172), .A3 (
           nx25181)) ;
    aoi22 ix25154 (.Y (nx25153), .A0 (camera_module_cache_ram_2__4), .A1 (
          nx35814), .B0 (camera_module_cache_ram_18__4), .B1 (nx35854)) ;
    dffr camera_module_cache_reg_ram_2__4 (.Q (camera_module_cache_ram_2__4), .QB (
         \$dummy [316]), .D (nx13773), .CLK (clk), .R (rst)) ;
    mux21_ni ix13774 (.Y (nx13773), .A0 (camera_module_cache_ram_2__4), .A1 (
             nx35376), .S0 (nx34994)) ;
    dffr camera_module_cache_reg_ram_18__4 (.Q (camera_module_cache_ram_18__4), 
         .QB (\$dummy [317]), .D (nx13763), .CLK (clk), .R (rst)) ;
    mux21_ni ix13764 (.Y (nx13763), .A0 (camera_module_cache_ram_18__4), .A1 (
             nx35376), .S0 (nx34990)) ;
    aoi22 ix25163 (.Y (nx25162), .A0 (camera_module_cache_ram_34__4), .A1 (
          nx35894), .B0 (camera_module_cache_ram_50__4), .B1 (nx35934)) ;
    dffr camera_module_cache_reg_ram_34__4 (.Q (camera_module_cache_ram_34__4), 
         .QB (\$dummy [318]), .D (nx13753), .CLK (clk), .R (rst)) ;
    mux21_ni ix13754 (.Y (nx13753), .A0 (camera_module_cache_ram_34__4), .A1 (
             nx35376), .S0 (nx34986)) ;
    dffr camera_module_cache_reg_ram_50__4 (.Q (camera_module_cache_ram_50__4), 
         .QB (\$dummy [319]), .D (nx13743), .CLK (clk), .R (rst)) ;
    mux21_ni ix13744 (.Y (nx13743), .A0 (camera_module_cache_ram_50__4), .A1 (
             nx35378), .S0 (nx34982)) ;
    aoi22 ix25173 (.Y (nx25172), .A0 (camera_module_cache_ram_66__4), .A1 (
          nx35974), .B0 (camera_module_cache_ram_82__4), .B1 (nx36014)) ;
    dffr camera_module_cache_reg_ram_66__4 (.Q (camera_module_cache_ram_66__4), 
         .QB (\$dummy [320]), .D (nx13733), .CLK (clk), .R (rst)) ;
    mux21_ni ix13734 (.Y (nx13733), .A0 (camera_module_cache_ram_66__4), .A1 (
             nx35378), .S0 (nx34978)) ;
    dffr camera_module_cache_reg_ram_82__4 (.Q (camera_module_cache_ram_82__4), 
         .QB (\$dummy [321]), .D (nx13723), .CLK (clk), .R (rst)) ;
    mux21_ni ix13724 (.Y (nx13723), .A0 (camera_module_cache_ram_82__4), .A1 (
             nx35378), .S0 (nx34974)) ;
    aoi22 ix25182 (.Y (nx25181), .A0 (camera_module_cache_ram_114__4), .A1 (
          nx36054), .B0 (camera_module_cache_ram_98__4), .B1 (nx36094)) ;
    dffr camera_module_cache_reg_ram_114__4 (.Q (camera_module_cache_ram_114__4)
         , .QB (\$dummy [322]), .D (nx13703), .CLK (clk), .R (rst)) ;
    mux21_ni ix13704 (.Y (nx13703), .A0 (camera_module_cache_ram_114__4), .A1 (
             nx35378), .S0 (nx34966)) ;
    dffr camera_module_cache_reg_ram_98__4 (.Q (camera_module_cache_ram_98__4), 
         .QB (\$dummy [323]), .D (nx13713), .CLK (clk), .R (rst)) ;
    mux21_ni ix13714 (.Y (nx13713), .A0 (camera_module_cache_ram_98__4), .A1 (
             nx35378), .S0 (nx34970)) ;
    nand04 ix16627 (.Y (nx16626), .A0 (nx25191), .A1 (nx25201), .A2 (nx25209), .A3 (
           nx25218)) ;
    aoi22 ix25192 (.Y (nx25191), .A0 (camera_module_cache_ram_130__4), .A1 (
          nx36134), .B0 (camera_module_cache_ram_146__4), .B1 (nx36174)) ;
    dffr camera_module_cache_reg_ram_130__4 (.Q (camera_module_cache_ram_130__4)
         , .QB (\$dummy [324]), .D (nx13693), .CLK (clk), .R (rst)) ;
    mux21_ni ix13694 (.Y (nx13693), .A0 (camera_module_cache_ram_130__4), .A1 (
             nx35378), .S0 (nx34962)) ;
    dffr camera_module_cache_reg_ram_146__4 (.Q (camera_module_cache_ram_146__4)
         , .QB (\$dummy [325]), .D (nx13683), .CLK (clk), .R (rst)) ;
    mux21_ni ix13684 (.Y (nx13683), .A0 (camera_module_cache_ram_146__4), .A1 (
             nx35378), .S0 (nx34958)) ;
    aoi22 ix25202 (.Y (nx25201), .A0 (camera_module_cache_ram_178__4), .A1 (
          nx36214), .B0 (camera_module_cache_ram_162__4), .B1 (nx36254)) ;
    dffr camera_module_cache_reg_ram_178__4 (.Q (camera_module_cache_ram_178__4)
         , .QB (\$dummy [326]), .D (nx13663), .CLK (clk), .R (rst)) ;
    mux21_ni ix13664 (.Y (nx13663), .A0 (camera_module_cache_ram_178__4), .A1 (
             nx35380), .S0 (nx34950)) ;
    dffr camera_module_cache_reg_ram_162__4 (.Q (camera_module_cache_ram_162__4)
         , .QB (\$dummy [327]), .D (nx13673), .CLK (clk), .R (rst)) ;
    mux21_ni ix13674 (.Y (nx13673), .A0 (camera_module_cache_ram_162__4), .A1 (
             nx35380), .S0 (nx34954)) ;
    aoi22 ix25210 (.Y (nx25209), .A0 (camera_module_cache_ram_194__4), .A1 (
          nx36294), .B0 (camera_module_cache_ram_210__4), .B1 (nx36334)) ;
    dffr camera_module_cache_reg_ram_194__4 (.Q (camera_module_cache_ram_194__4)
         , .QB (\$dummy [328]), .D (nx13653), .CLK (clk), .R (rst)) ;
    mux21_ni ix13654 (.Y (nx13653), .A0 (camera_module_cache_ram_194__4), .A1 (
             nx35380), .S0 (nx34946)) ;
    dffr camera_module_cache_reg_ram_210__4 (.Q (camera_module_cache_ram_210__4)
         , .QB (\$dummy [329]), .D (nx13643), .CLK (clk), .R (rst)) ;
    mux21_ni ix13644 (.Y (nx13643), .A0 (camera_module_cache_ram_210__4), .A1 (
             nx35380), .S0 (nx34942)) ;
    aoi22 ix25219 (.Y (nx25218), .A0 (camera_module_cache_ram_226__4), .A1 (
          nx36374), .B0 (camera_module_cache_ram_242__4), .B1 (nx36414)) ;
    dffr camera_module_cache_reg_ram_226__4 (.Q (camera_module_cache_ram_226__4)
         , .QB (\$dummy [330]), .D (nx13633), .CLK (clk), .R (rst)) ;
    mux21_ni ix13634 (.Y (nx13633), .A0 (camera_module_cache_ram_226__4), .A1 (
             nx35380), .S0 (nx34938)) ;
    dffr camera_module_cache_reg_ram_242__4 (.Q (camera_module_cache_ram_242__4)
         , .QB (\$dummy [331]), .D (nx13623), .CLK (clk), .R (rst)) ;
    mux21_ni ix13624 (.Y (nx13623), .A0 (camera_module_cache_ram_242__4), .A1 (
             nx35380), .S0 (nx34934)) ;
    oai21 ix25228 (.Y (nx25227), .A0 (nx16542), .A1 (nx16464), .B0 (nx36460)) ;
    nand04 ix16543 (.Y (nx16542), .A0 (nx25231), .A1 (nx25241), .A2 (nx25251), .A3 (
           nx25261)) ;
    aoi22 ix25232 (.Y (nx25231), .A0 (camera_module_cache_ram_3__4), .A1 (
          nx35814), .B0 (camera_module_cache_ram_19__4), .B1 (nx35854)) ;
    dffr camera_module_cache_reg_ram_3__4 (.Q (camera_module_cache_ram_3__4), .QB (
         \$dummy [332]), .D (nx13613), .CLK (clk), .R (rst)) ;
    mux21_ni ix13614 (.Y (nx13613), .A0 (camera_module_cache_ram_3__4), .A1 (
             nx35380), .S0 (nx34924)) ;
    dffr camera_module_cache_reg_ram_19__4 (.Q (camera_module_cache_ram_19__4), 
         .QB (\$dummy [333]), .D (nx13603), .CLK (clk), .R (rst)) ;
    mux21_ni ix13604 (.Y (nx13603), .A0 (camera_module_cache_ram_19__4), .A1 (
             nx35382), .S0 (nx34920)) ;
    aoi22 ix25242 (.Y (nx25241), .A0 (camera_module_cache_ram_35__4), .A1 (
          nx35894), .B0 (camera_module_cache_ram_51__4), .B1 (nx35934)) ;
    dffr camera_module_cache_reg_ram_35__4 (.Q (camera_module_cache_ram_35__4), 
         .QB (\$dummy [334]), .D (nx13593), .CLK (clk), .R (rst)) ;
    mux21_ni ix13594 (.Y (nx13593), .A0 (camera_module_cache_ram_35__4), .A1 (
             nx35382), .S0 (nx34916)) ;
    dffr camera_module_cache_reg_ram_51__4 (.Q (camera_module_cache_ram_51__4), 
         .QB (\$dummy [335]), .D (nx13583), .CLK (clk), .R (rst)) ;
    mux21_ni ix13584 (.Y (nx13583), .A0 (camera_module_cache_ram_51__4), .A1 (
             nx35382), .S0 (nx34912)) ;
    aoi22 ix25252 (.Y (nx25251), .A0 (camera_module_cache_ram_67__4), .A1 (
          nx35974), .B0 (camera_module_cache_ram_83__4), .B1 (nx36014)) ;
    dffr camera_module_cache_reg_ram_67__4 (.Q (camera_module_cache_ram_67__4), 
         .QB (\$dummy [336]), .D (nx13573), .CLK (clk), .R (rst)) ;
    mux21_ni ix13574 (.Y (nx13573), .A0 (camera_module_cache_ram_67__4), .A1 (
             nx35382), .S0 (nx34908)) ;
    dffr camera_module_cache_reg_ram_83__4 (.Q (camera_module_cache_ram_83__4), 
         .QB (\$dummy [337]), .D (nx13563), .CLK (clk), .R (rst)) ;
    mux21_ni ix13564 (.Y (nx13563), .A0 (camera_module_cache_ram_83__4), .A1 (
             nx35382), .S0 (nx34904)) ;
    aoi22 ix25262 (.Y (nx25261), .A0 (camera_module_cache_ram_115__4), .A1 (
          nx36054), .B0 (camera_module_cache_ram_99__4), .B1 (nx36094)) ;
    dffr camera_module_cache_reg_ram_115__4 (.Q (camera_module_cache_ram_115__4)
         , .QB (\$dummy [338]), .D (nx13543), .CLK (clk), .R (rst)) ;
    mux21_ni ix13544 (.Y (nx13543), .A0 (camera_module_cache_ram_115__4), .A1 (
             nx35382), .S0 (nx34896)) ;
    dffr camera_module_cache_reg_ram_99__4 (.Q (camera_module_cache_ram_99__4), 
         .QB (\$dummy [339]), .D (nx13553), .CLK (clk), .R (rst)) ;
    mux21_ni ix13554 (.Y (nx13553), .A0 (camera_module_cache_ram_99__4), .A1 (
             nx35382), .S0 (nx34900)) ;
    nand04 ix16465 (.Y (nx16464), .A0 (nx25271), .A1 (nx25281), .A2 (nx25291), .A3 (
           nx25301)) ;
    aoi22 ix25272 (.Y (nx25271), .A0 (camera_module_cache_ram_131__4), .A1 (
          nx36134), .B0 (camera_module_cache_ram_147__4), .B1 (nx36174)) ;
    dffr camera_module_cache_reg_ram_131__4 (.Q (camera_module_cache_ram_131__4)
         , .QB (\$dummy [340]), .D (nx13533), .CLK (clk), .R (rst)) ;
    mux21_ni ix13534 (.Y (nx13533), .A0 (camera_module_cache_ram_131__4), .A1 (
             nx35384), .S0 (nx34892)) ;
    dffr camera_module_cache_reg_ram_147__4 (.Q (camera_module_cache_ram_147__4)
         , .QB (\$dummy [341]), .D (nx13523), .CLK (clk), .R (rst)) ;
    mux21_ni ix13524 (.Y (nx13523), .A0 (camera_module_cache_ram_147__4), .A1 (
             nx35384), .S0 (nx34888)) ;
    aoi22 ix25282 (.Y (nx25281), .A0 (camera_module_cache_ram_179__4), .A1 (
          nx36214), .B0 (camera_module_cache_ram_163__4), .B1 (nx36254)) ;
    dffr camera_module_cache_reg_ram_179__4 (.Q (camera_module_cache_ram_179__4)
         , .QB (\$dummy [342]), .D (nx13503), .CLK (clk), .R (rst)) ;
    mux21_ni ix13504 (.Y (nx13503), .A0 (camera_module_cache_ram_179__4), .A1 (
             nx35384), .S0 (nx34880)) ;
    dffr camera_module_cache_reg_ram_163__4 (.Q (camera_module_cache_ram_163__4)
         , .QB (\$dummy [343]), .D (nx13513), .CLK (clk), .R (rst)) ;
    mux21_ni ix13514 (.Y (nx13513), .A0 (camera_module_cache_ram_163__4), .A1 (
             nx35384), .S0 (nx34884)) ;
    aoi22 ix25292 (.Y (nx25291), .A0 (camera_module_cache_ram_195__4), .A1 (
          nx36294), .B0 (camera_module_cache_ram_211__4), .B1 (nx36334)) ;
    dffr camera_module_cache_reg_ram_195__4 (.Q (camera_module_cache_ram_195__4)
         , .QB (\$dummy [344]), .D (nx13493), .CLK (clk), .R (rst)) ;
    mux21_ni ix13494 (.Y (nx13493), .A0 (camera_module_cache_ram_195__4), .A1 (
             nx35384), .S0 (nx34876)) ;
    dffr camera_module_cache_reg_ram_211__4 (.Q (camera_module_cache_ram_211__4)
         , .QB (\$dummy [345]), .D (nx13483), .CLK (clk), .R (rst)) ;
    mux21_ni ix13484 (.Y (nx13483), .A0 (camera_module_cache_ram_211__4), .A1 (
             nx35384), .S0 (nx34872)) ;
    aoi22 ix25302 (.Y (nx25301), .A0 (camera_module_cache_ram_227__4), .A1 (
          nx36374), .B0 (camera_module_cache_ram_243__4), .B1 (nx36414)) ;
    dffr camera_module_cache_reg_ram_227__4 (.Q (camera_module_cache_ram_227__4)
         , .QB (\$dummy [346]), .D (nx13473), .CLK (clk), .R (rst)) ;
    mux21_ni ix13474 (.Y (nx13473), .A0 (camera_module_cache_ram_227__4), .A1 (
             nx35384), .S0 (nx34868)) ;
    dffr camera_module_cache_reg_ram_243__4 (.Q (camera_module_cache_ram_243__4)
         , .QB (\$dummy [347]), .D (nx13463), .CLK (clk), .R (rst)) ;
    mux21_ni ix13464 (.Y (nx13463), .A0 (camera_module_cache_ram_243__4), .A1 (
             nx35386), .S0 (nx34864)) ;
    nand04 ix16387 (.Y (nx16386), .A0 (nx25311), .A1 (nx25397), .A2 (nx25489), .A3 (
           nx25576)) ;
    oai21 ix25312 (.Y (nx25311), .A0 (nx16376), .A1 (nx16298), .B0 (nx36464)) ;
    nand04 ix16377 (.Y (nx16376), .A0 (nx25315), .A1 (nx25324), .A2 (nx25334), .A3 (
           nx25343)) ;
    aoi22 ix25316 (.Y (nx25315), .A0 (camera_module_cache_ram_4__4), .A1 (
          nx35814), .B0 (camera_module_cache_ram_20__4), .B1 (nx35854)) ;
    dffr camera_module_cache_reg_ram_4__4 (.Q (camera_module_cache_ram_4__4), .QB (
         \$dummy [348]), .D (nx13453), .CLK (clk), .R (rst)) ;
    mux21_ni ix13454 (.Y (nx13453), .A0 (camera_module_cache_ram_4__4), .A1 (
             nx35386), .S0 (nx34854)) ;
    dffr camera_module_cache_reg_ram_20__4 (.Q (camera_module_cache_ram_20__4), 
         .QB (\$dummy [349]), .D (nx13443), .CLK (clk), .R (rst)) ;
    mux21_ni ix13444 (.Y (nx13443), .A0 (camera_module_cache_ram_20__4), .A1 (
             nx35386), .S0 (nx34850)) ;
    aoi22 ix25325 (.Y (nx25324), .A0 (camera_module_cache_ram_36__4), .A1 (
          nx35894), .B0 (camera_module_cache_ram_52__4), .B1 (nx35934)) ;
    dffr camera_module_cache_reg_ram_36__4 (.Q (camera_module_cache_ram_36__4), 
         .QB (\$dummy [350]), .D (nx13433), .CLK (clk), .R (rst)) ;
    mux21_ni ix13434 (.Y (nx13433), .A0 (camera_module_cache_ram_36__4), .A1 (
             nx35386), .S0 (nx34846)) ;
    dffr camera_module_cache_reg_ram_52__4 (.Q (camera_module_cache_ram_52__4), 
         .QB (\$dummy [351]), .D (nx13423), .CLK (clk), .R (rst)) ;
    mux21_ni ix13424 (.Y (nx13423), .A0 (camera_module_cache_ram_52__4), .A1 (
             nx35386), .S0 (nx34842)) ;
    aoi22 ix25335 (.Y (nx25334), .A0 (camera_module_cache_ram_68__4), .A1 (
          nx35974), .B0 (camera_module_cache_ram_84__4), .B1 (nx36014)) ;
    dffr camera_module_cache_reg_ram_68__4 (.Q (camera_module_cache_ram_68__4), 
         .QB (\$dummy [352]), .D (nx13413), .CLK (clk), .R (rst)) ;
    mux21_ni ix13414 (.Y (nx13413), .A0 (camera_module_cache_ram_68__4), .A1 (
             nx35386), .S0 (nx34838)) ;
    dffr camera_module_cache_reg_ram_84__4 (.Q (camera_module_cache_ram_84__4), 
         .QB (\$dummy [353]), .D (nx13403), .CLK (clk), .R (rst)) ;
    mux21_ni ix13404 (.Y (nx13403), .A0 (camera_module_cache_ram_84__4), .A1 (
             nx35386), .S0 (nx34834)) ;
    aoi22 ix25344 (.Y (nx25343), .A0 (camera_module_cache_ram_116__4), .A1 (
          nx36054), .B0 (camera_module_cache_ram_100__4), .B1 (nx36094)) ;
    dffr camera_module_cache_reg_ram_116__4 (.Q (camera_module_cache_ram_116__4)
         , .QB (\$dummy [354]), .D (nx13383), .CLK (clk), .R (rst)) ;
    mux21_ni ix13384 (.Y (nx13383), .A0 (camera_module_cache_ram_116__4), .A1 (
             nx35388), .S0 (nx34826)) ;
    dffr camera_module_cache_reg_ram_100__4 (.Q (camera_module_cache_ram_100__4)
         , .QB (\$dummy [355]), .D (nx13393), .CLK (clk), .R (rst)) ;
    mux21_ni ix13394 (.Y (nx13393), .A0 (camera_module_cache_ram_100__4), .A1 (
             nx35388), .S0 (nx34830)) ;
    nand04 ix16299 (.Y (nx16298), .A0 (nx25353), .A1 (nx25365), .A2 (nx25376), .A3 (
           nx25386)) ;
    aoi22 ix25354 (.Y (nx25353), .A0 (camera_module_cache_ram_132__4), .A1 (
          nx36134), .B0 (camera_module_cache_ram_148__4), .B1 (nx36174)) ;
    dffr camera_module_cache_reg_ram_132__4 (.Q (camera_module_cache_ram_132__4)
         , .QB (\$dummy [356]), .D (nx13373), .CLK (clk), .R (rst)) ;
    mux21_ni ix13374 (.Y (nx13373), .A0 (camera_module_cache_ram_132__4), .A1 (
             nx35388), .S0 (nx34822)) ;
    dffr camera_module_cache_reg_ram_148__4 (.Q (camera_module_cache_ram_148__4)
         , .QB (\$dummy [357]), .D (nx13363), .CLK (clk), .R (rst)) ;
    mux21_ni ix13364 (.Y (nx13363), .A0 (camera_module_cache_ram_148__4), .A1 (
             nx35388), .S0 (nx34818)) ;
    aoi22 ix25366 (.Y (nx25365), .A0 (camera_module_cache_ram_180__4), .A1 (
          nx36214), .B0 (camera_module_cache_ram_164__4), .B1 (nx36254)) ;
    dffr camera_module_cache_reg_ram_180__4 (.Q (camera_module_cache_ram_180__4)
         , .QB (\$dummy [358]), .D (nx13343), .CLK (clk), .R (rst)) ;
    mux21_ni ix13344 (.Y (nx13343), .A0 (camera_module_cache_ram_180__4), .A1 (
             nx35388), .S0 (nx34810)) ;
    dffr camera_module_cache_reg_ram_164__4 (.Q (camera_module_cache_ram_164__4)
         , .QB (\$dummy [359]), .D (nx13353), .CLK (clk), .R (rst)) ;
    mux21_ni ix13354 (.Y (nx13353), .A0 (camera_module_cache_ram_164__4), .A1 (
             nx35388), .S0 (nx34814)) ;
    aoi22 ix25377 (.Y (nx25376), .A0 (camera_module_cache_ram_196__4), .A1 (
          nx36294), .B0 (camera_module_cache_ram_212__4), .B1 (nx36334)) ;
    dffr camera_module_cache_reg_ram_196__4 (.Q (camera_module_cache_ram_196__4)
         , .QB (\$dummy [360]), .D (nx13333), .CLK (clk), .R (rst)) ;
    mux21_ni ix13334 (.Y (nx13333), .A0 (camera_module_cache_ram_196__4), .A1 (
             nx35388), .S0 (nx34806)) ;
    dffr camera_module_cache_reg_ram_212__4 (.Q (camera_module_cache_ram_212__4)
         , .QB (\$dummy [361]), .D (nx13323), .CLK (clk), .R (rst)) ;
    mux21_ni ix13324 (.Y (nx13323), .A0 (camera_module_cache_ram_212__4), .A1 (
             nx35390), .S0 (nx34802)) ;
    aoi22 ix25387 (.Y (nx25386), .A0 (camera_module_cache_ram_228__4), .A1 (
          nx36374), .B0 (camera_module_cache_ram_244__4), .B1 (nx36414)) ;
    dffr camera_module_cache_reg_ram_228__4 (.Q (camera_module_cache_ram_228__4)
         , .QB (\$dummy [362]), .D (nx13313), .CLK (clk), .R (rst)) ;
    mux21_ni ix13314 (.Y (nx13313), .A0 (camera_module_cache_ram_228__4), .A1 (
             nx35390), .S0 (nx34798)) ;
    dffr camera_module_cache_reg_ram_244__4 (.Q (camera_module_cache_ram_244__4)
         , .QB (\$dummy [363]), .D (nx13303), .CLK (clk), .R (rst)) ;
    mux21_ni ix13304 (.Y (nx13303), .A0 (camera_module_cache_ram_244__4), .A1 (
             nx35390), .S0 (nx34794)) ;
    oai21 ix25398 (.Y (nx25397), .A0 (nx16214), .A1 (nx16136), .B0 (nx36468)) ;
    nand04 ix16215 (.Y (nx16214), .A0 (nx25401), .A1 (nx25413), .A2 (nx25425), .A3 (
           nx25437)) ;
    aoi22 ix25402 (.Y (nx25401), .A0 (camera_module_cache_ram_5__4), .A1 (
          nx35814), .B0 (camera_module_cache_ram_21__4), .B1 (nx35854)) ;
    dffr camera_module_cache_reg_ram_5__4 (.Q (camera_module_cache_ram_5__4), .QB (
         \$dummy [364]), .D (nx13293), .CLK (clk), .R (rst)) ;
    mux21_ni ix13294 (.Y (nx13293), .A0 (camera_module_cache_ram_5__4), .A1 (
             nx35390), .S0 (nx34784)) ;
    dffr camera_module_cache_reg_ram_21__4 (.Q (camera_module_cache_ram_21__4), 
         .QB (\$dummy [365]), .D (nx13283), .CLK (clk), .R (rst)) ;
    mux21_ni ix13284 (.Y (nx13283), .A0 (camera_module_cache_ram_21__4), .A1 (
             nx35390), .S0 (nx34780)) ;
    aoi22 ix25414 (.Y (nx25413), .A0 (camera_module_cache_ram_37__4), .A1 (
          nx35894), .B0 (camera_module_cache_ram_53__4), .B1 (nx35934)) ;
    dffr camera_module_cache_reg_ram_37__4 (.Q (camera_module_cache_ram_37__4), 
         .QB (\$dummy [366]), .D (nx13273), .CLK (clk), .R (rst)) ;
    mux21_ni ix13274 (.Y (nx13273), .A0 (camera_module_cache_ram_37__4), .A1 (
             nx35390), .S0 (nx34776)) ;
    dffr camera_module_cache_reg_ram_53__4 (.Q (camera_module_cache_ram_53__4), 
         .QB (\$dummy [367]), .D (nx13263), .CLK (clk), .R (rst)) ;
    mux21_ni ix13264 (.Y (nx13263), .A0 (camera_module_cache_ram_53__4), .A1 (
             nx35390), .S0 (nx34772)) ;
    aoi22 ix25426 (.Y (nx25425), .A0 (camera_module_cache_ram_69__4), .A1 (
          nx35974), .B0 (camera_module_cache_ram_85__4), .B1 (nx36014)) ;
    dffr camera_module_cache_reg_ram_69__4 (.Q (camera_module_cache_ram_69__4), 
         .QB (\$dummy [368]), .D (nx13253), .CLK (clk), .R (rst)) ;
    mux21_ni ix13254 (.Y (nx13253), .A0 (camera_module_cache_ram_69__4), .A1 (
             nx35392), .S0 (nx34768)) ;
    dffr camera_module_cache_reg_ram_85__4 (.Q (camera_module_cache_ram_85__4), 
         .QB (\$dummy [369]), .D (nx13243), .CLK (clk), .R (rst)) ;
    mux21_ni ix13244 (.Y (nx13243), .A0 (camera_module_cache_ram_85__4), .A1 (
             nx35392), .S0 (nx34764)) ;
    aoi22 ix25438 (.Y (nx25437), .A0 (camera_module_cache_ram_117__4), .A1 (
          nx36054), .B0 (camera_module_cache_ram_101__4), .B1 (nx36094)) ;
    dffr camera_module_cache_reg_ram_117__4 (.Q (camera_module_cache_ram_117__4)
         , .QB (\$dummy [370]), .D (nx13223), .CLK (clk), .R (rst)) ;
    mux21_ni ix13224 (.Y (nx13223), .A0 (camera_module_cache_ram_117__4), .A1 (
             nx35392), .S0 (nx34756)) ;
    dffr camera_module_cache_reg_ram_101__4 (.Q (camera_module_cache_ram_101__4)
         , .QB (\$dummy [371]), .D (nx13233), .CLK (clk), .R (rst)) ;
    mux21_ni ix13234 (.Y (nx13233), .A0 (camera_module_cache_ram_101__4), .A1 (
             nx35392), .S0 (nx34760)) ;
    nand04 ix16137 (.Y (nx16136), .A0 (nx25449), .A1 (nx25459), .A2 (nx25469), .A3 (
           nx25480)) ;
    aoi22 ix25450 (.Y (nx25449), .A0 (camera_module_cache_ram_133__4), .A1 (
          nx36134), .B0 (camera_module_cache_ram_149__4), .B1 (nx36174)) ;
    dffr camera_module_cache_reg_ram_133__4 (.Q (camera_module_cache_ram_133__4)
         , .QB (\$dummy [372]), .D (nx13213), .CLK (clk), .R (rst)) ;
    mux21_ni ix13214 (.Y (nx13213), .A0 (camera_module_cache_ram_133__4), .A1 (
             nx35392), .S0 (nx34752)) ;
    dffr camera_module_cache_reg_ram_149__4 (.Q (camera_module_cache_ram_149__4)
         , .QB (\$dummy [373]), .D (nx13203), .CLK (clk), .R (rst)) ;
    mux21_ni ix13204 (.Y (nx13203), .A0 (camera_module_cache_ram_149__4), .A1 (
             nx35392), .S0 (nx34748)) ;
    aoi22 ix25460 (.Y (nx25459), .A0 (camera_module_cache_ram_181__4), .A1 (
          nx36214), .B0 (camera_module_cache_ram_165__4), .B1 (nx36254)) ;
    dffr camera_module_cache_reg_ram_181__4 (.Q (camera_module_cache_ram_181__4)
         , .QB (\$dummy [374]), .D (nx13183), .CLK (clk), .R (rst)) ;
    mux21_ni ix13184 (.Y (nx13183), .A0 (camera_module_cache_ram_181__4), .A1 (
             nx35392), .S0 (nx34740)) ;
    dffr camera_module_cache_reg_ram_165__4 (.Q (camera_module_cache_ram_165__4)
         , .QB (\$dummy [375]), .D (nx13193), .CLK (clk), .R (rst)) ;
    mux21_ni ix13194 (.Y (nx13193), .A0 (camera_module_cache_ram_165__4), .A1 (
             nx35394), .S0 (nx34744)) ;
    aoi22 ix25470 (.Y (nx25469), .A0 (camera_module_cache_ram_197__4), .A1 (
          nx36294), .B0 (camera_module_cache_ram_213__4), .B1 (nx36334)) ;
    dffr camera_module_cache_reg_ram_197__4 (.Q (camera_module_cache_ram_197__4)
         , .QB (\$dummy [376]), .D (nx13173), .CLK (clk), .R (rst)) ;
    mux21_ni ix13174 (.Y (nx13173), .A0 (camera_module_cache_ram_197__4), .A1 (
             nx35394), .S0 (nx34736)) ;
    dffr camera_module_cache_reg_ram_213__4 (.Q (camera_module_cache_ram_213__4)
         , .QB (\$dummy [377]), .D (nx13163), .CLK (clk), .R (rst)) ;
    mux21_ni ix13164 (.Y (nx13163), .A0 (camera_module_cache_ram_213__4), .A1 (
             nx35394), .S0 (nx34732)) ;
    aoi22 ix25481 (.Y (nx25480), .A0 (camera_module_cache_ram_229__4), .A1 (
          nx36374), .B0 (camera_module_cache_ram_245__4), .B1 (nx36414)) ;
    dffr camera_module_cache_reg_ram_229__4 (.Q (camera_module_cache_ram_229__4)
         , .QB (\$dummy [378]), .D (nx13153), .CLK (clk), .R (rst)) ;
    mux21_ni ix13154 (.Y (nx13153), .A0 (camera_module_cache_ram_229__4), .A1 (
             nx35394), .S0 (nx34728)) ;
    dffr camera_module_cache_reg_ram_245__4 (.Q (camera_module_cache_ram_245__4)
         , .QB (\$dummy [379]), .D (nx13143), .CLK (clk), .R (rst)) ;
    mux21_ni ix13144 (.Y (nx13143), .A0 (camera_module_cache_ram_245__4), .A1 (
             nx35394), .S0 (nx34724)) ;
    oai21 ix25490 (.Y (nx25489), .A0 (nx16050), .A1 (nx15972), .B0 (nx36472)) ;
    nand04 ix16051 (.Y (nx16050), .A0 (nx25493), .A1 (nx25502), .A2 (nx25515), .A3 (
           nx25525)) ;
    aoi22 ix25494 (.Y (nx25493), .A0 (camera_module_cache_ram_6__4), .A1 (
          nx35814), .B0 (camera_module_cache_ram_22__4), .B1 (nx35854)) ;
    dffr camera_module_cache_reg_ram_6__4 (.Q (camera_module_cache_ram_6__4), .QB (
         \$dummy [380]), .D (nx13133), .CLK (clk), .R (rst)) ;
    mux21_ni ix13134 (.Y (nx13133), .A0 (camera_module_cache_ram_6__4), .A1 (
             nx35394), .S0 (nx34714)) ;
    dffr camera_module_cache_reg_ram_22__4 (.Q (camera_module_cache_ram_22__4), 
         .QB (\$dummy [381]), .D (nx13123), .CLK (clk), .R (rst)) ;
    mux21_ni ix13124 (.Y (nx13123), .A0 (camera_module_cache_ram_22__4), .A1 (
             nx35394), .S0 (nx34710)) ;
    aoi22 ix25504 (.Y (nx25502), .A0 (camera_module_cache_ram_38__4), .A1 (
          nx35894), .B0 (camera_module_cache_ram_54__4), .B1 (nx35934)) ;
    dffr camera_module_cache_reg_ram_38__4 (.Q (camera_module_cache_ram_38__4), 
         .QB (\$dummy [382]), .D (nx13113), .CLK (clk), .R (rst)) ;
    mux21_ni ix13114 (.Y (nx13113), .A0 (camera_module_cache_ram_38__4), .A1 (
             nx35396), .S0 (nx34706)) ;
    dffr camera_module_cache_reg_ram_54__4 (.Q (camera_module_cache_ram_54__4), 
         .QB (\$dummy [383]), .D (nx13103), .CLK (clk), .R (rst)) ;
    mux21_ni ix13104 (.Y (nx13103), .A0 (camera_module_cache_ram_54__4), .A1 (
             nx35396), .S0 (nx34702)) ;
    aoi22 ix25516 (.Y (nx25515), .A0 (camera_module_cache_ram_70__4), .A1 (
          nx35974), .B0 (camera_module_cache_ram_86__4), .B1 (nx36014)) ;
    dffr camera_module_cache_reg_ram_70__4 (.Q (camera_module_cache_ram_70__4), 
         .QB (\$dummy [384]), .D (nx13093), .CLK (clk), .R (rst)) ;
    mux21_ni ix13094 (.Y (nx13093), .A0 (camera_module_cache_ram_70__4), .A1 (
             nx35396), .S0 (nx34698)) ;
    dffr camera_module_cache_reg_ram_86__4 (.Q (camera_module_cache_ram_86__4), 
         .QB (\$dummy [385]), .D (nx13083), .CLK (clk), .R (rst)) ;
    mux21_ni ix13084 (.Y (nx13083), .A0 (camera_module_cache_ram_86__4), .A1 (
             nx35396), .S0 (nx34694)) ;
    aoi22 ix25526 (.Y (nx25525), .A0 (camera_module_cache_ram_118__4), .A1 (
          nx36054), .B0 (camera_module_cache_ram_102__4), .B1 (nx36094)) ;
    dffr camera_module_cache_reg_ram_118__4 (.Q (camera_module_cache_ram_118__4)
         , .QB (\$dummy [386]), .D (nx13063), .CLK (clk), .R (rst)) ;
    mux21_ni ix13064 (.Y (nx13063), .A0 (camera_module_cache_ram_118__4), .A1 (
             nx35396), .S0 (nx34686)) ;
    dffr camera_module_cache_reg_ram_102__4 (.Q (camera_module_cache_ram_102__4)
         , .QB (\$dummy [387]), .D (nx13073), .CLK (clk), .R (rst)) ;
    mux21_ni ix13074 (.Y (nx13073), .A0 (camera_module_cache_ram_102__4), .A1 (
             nx35396), .S0 (nx34690)) ;
    nand04 ix15973 (.Y (nx15972), .A0 (nx25536), .A1 (nx25549), .A2 (nx25559), .A3 (
           nx25568)) ;
    aoi22 ix25538 (.Y (nx25536), .A0 (camera_module_cache_ram_134__4), .A1 (
          nx36134), .B0 (camera_module_cache_ram_150__4), .B1 (nx36174)) ;
    dffr camera_module_cache_reg_ram_134__4 (.Q (camera_module_cache_ram_134__4)
         , .QB (\$dummy [388]), .D (nx13053), .CLK (clk), .R (rst)) ;
    mux21_ni ix13054 (.Y (nx13053), .A0 (camera_module_cache_ram_134__4), .A1 (
             nx35396), .S0 (nx34682)) ;
    dffr camera_module_cache_reg_ram_150__4 (.Q (camera_module_cache_ram_150__4)
         , .QB (\$dummy [389]), .D (nx13043), .CLK (clk), .R (rst)) ;
    mux21_ni ix13044 (.Y (nx13043), .A0 (camera_module_cache_ram_150__4), .A1 (
             nx35398), .S0 (nx34678)) ;
    aoi22 ix25550 (.Y (nx25549), .A0 (camera_module_cache_ram_182__4), .A1 (
          nx36214), .B0 (camera_module_cache_ram_166__4), .B1 (nx36254)) ;
    dffr camera_module_cache_reg_ram_182__4 (.Q (camera_module_cache_ram_182__4)
         , .QB (\$dummy [390]), .D (nx13023), .CLK (clk), .R (rst)) ;
    mux21_ni ix13024 (.Y (nx13023), .A0 (camera_module_cache_ram_182__4), .A1 (
             nx35398), .S0 (nx34670)) ;
    dffr camera_module_cache_reg_ram_166__4 (.Q (camera_module_cache_ram_166__4)
         , .QB (\$dummy [391]), .D (nx13033), .CLK (clk), .R (rst)) ;
    mux21_ni ix13034 (.Y (nx13033), .A0 (camera_module_cache_ram_166__4), .A1 (
             nx35398), .S0 (nx34674)) ;
    aoi22 ix25560 (.Y (nx25559), .A0 (camera_module_cache_ram_198__4), .A1 (
          nx36294), .B0 (camera_module_cache_ram_214__4), .B1 (nx36334)) ;
    dffr camera_module_cache_reg_ram_198__4 (.Q (camera_module_cache_ram_198__4)
         , .QB (\$dummy [392]), .D (nx13013), .CLK (clk), .R (rst)) ;
    mux21_ni ix13014 (.Y (nx13013), .A0 (camera_module_cache_ram_198__4), .A1 (
             nx35398), .S0 (nx34666)) ;
    dffr camera_module_cache_reg_ram_214__4 (.Q (camera_module_cache_ram_214__4)
         , .QB (\$dummy [393]), .D (nx13003), .CLK (clk), .R (rst)) ;
    mux21_ni ix13004 (.Y (nx13003), .A0 (camera_module_cache_ram_214__4), .A1 (
             nx35398), .S0 (nx34662)) ;
    aoi22 ix25569 (.Y (nx25568), .A0 (camera_module_cache_ram_230__4), .A1 (
          nx36374), .B0 (camera_module_cache_ram_246__4), .B1 (nx36414)) ;
    dffr camera_module_cache_reg_ram_230__4 (.Q (camera_module_cache_ram_230__4)
         , .QB (\$dummy [394]), .D (nx12993), .CLK (clk), .R (rst)) ;
    mux21_ni ix12994 (.Y (nx12993), .A0 (camera_module_cache_ram_230__4), .A1 (
             nx35398), .S0 (nx34658)) ;
    dffr camera_module_cache_reg_ram_246__4 (.Q (camera_module_cache_ram_246__4)
         , .QB (\$dummy [395]), .D (nx12983), .CLK (clk), .R (rst)) ;
    mux21_ni ix12984 (.Y (nx12983), .A0 (camera_module_cache_ram_246__4), .A1 (
             nx35398), .S0 (nx34654)) ;
    oai21 ix25578 (.Y (nx25576), .A0 (nx15888), .A1 (nx15810), .B0 (nx36476)) ;
    nand04 ix15889 (.Y (nx15888), .A0 (nx25581), .A1 (nx25593), .A2 (nx25604), .A3 (
           nx25613)) ;
    aoi22 ix25582 (.Y (nx25581), .A0 (camera_module_cache_ram_7__4), .A1 (
          nx35814), .B0 (camera_module_cache_ram_23__4), .B1 (nx35854)) ;
    dffr camera_module_cache_reg_ram_7__4 (.Q (camera_module_cache_ram_7__4), .QB (
         \$dummy [396]), .D (nx12973), .CLK (clk), .R (rst)) ;
    mux21_ni ix12974 (.Y (nx12973), .A0 (camera_module_cache_ram_7__4), .A1 (
             nx35400), .S0 (nx34644)) ;
    dffr camera_module_cache_reg_ram_23__4 (.Q (camera_module_cache_ram_23__4), 
         .QB (\$dummy [397]), .D (nx12963), .CLK (clk), .R (rst)) ;
    mux21_ni ix12964 (.Y (nx12963), .A0 (camera_module_cache_ram_23__4), .A1 (
             nx35400), .S0 (nx34640)) ;
    aoi22 ix25594 (.Y (nx25593), .A0 (camera_module_cache_ram_39__4), .A1 (
          nx35894), .B0 (camera_module_cache_ram_55__4), .B1 (nx35934)) ;
    dffr camera_module_cache_reg_ram_39__4 (.Q (camera_module_cache_ram_39__4), 
         .QB (\$dummy [398]), .D (nx12953), .CLK (clk), .R (rst)) ;
    mux21_ni ix12954 (.Y (nx12953), .A0 (camera_module_cache_ram_39__4), .A1 (
             nx35400), .S0 (nx34636)) ;
    dffr camera_module_cache_reg_ram_55__4 (.Q (camera_module_cache_ram_55__4), 
         .QB (\$dummy [399]), .D (nx12943), .CLK (clk), .R (rst)) ;
    mux21_ni ix12944 (.Y (nx12943), .A0 (camera_module_cache_ram_55__4), .A1 (
             nx35400), .S0 (nx34632)) ;
    aoi22 ix25605 (.Y (nx25604), .A0 (camera_module_cache_ram_71__4), .A1 (
          nx35974), .B0 (camera_module_cache_ram_87__4), .B1 (nx36014)) ;
    dffr camera_module_cache_reg_ram_71__4 (.Q (camera_module_cache_ram_71__4), 
         .QB (\$dummy [400]), .D (nx12933), .CLK (clk), .R (rst)) ;
    mux21_ni ix12934 (.Y (nx12933), .A0 (camera_module_cache_ram_71__4), .A1 (
             nx35400), .S0 (nx34628)) ;
    dffr camera_module_cache_reg_ram_87__4 (.Q (camera_module_cache_ram_87__4), 
         .QB (\$dummy [401]), .D (nx12923), .CLK (clk), .R (rst)) ;
    mux21_ni ix12924 (.Y (nx12923), .A0 (camera_module_cache_ram_87__4), .A1 (
             nx35400), .S0 (nx34624)) ;
    aoi22 ix25614 (.Y (nx25613), .A0 (camera_module_cache_ram_119__4), .A1 (
          nx36054), .B0 (camera_module_cache_ram_103__4), .B1 (nx36094)) ;
    dffr camera_module_cache_reg_ram_119__4 (.Q (camera_module_cache_ram_119__4)
         , .QB (\$dummy [402]), .D (nx12903), .CLK (clk), .R (rst)) ;
    mux21_ni ix12904 (.Y (nx12903), .A0 (camera_module_cache_ram_119__4), .A1 (
             nx35400), .S0 (nx34616)) ;
    dffr camera_module_cache_reg_ram_103__4 (.Q (camera_module_cache_ram_103__4)
         , .QB (\$dummy [403]), .D (nx12913), .CLK (clk), .R (rst)) ;
    mux21_ni ix12914 (.Y (nx12913), .A0 (camera_module_cache_ram_103__4), .A1 (
             nx35402), .S0 (nx34620)) ;
    nand04 ix15811 (.Y (nx15810), .A0 (nx25625), .A1 (nx25634), .A2 (nx25644), .A3 (
           nx25655)) ;
    aoi22 ix25626 (.Y (nx25625), .A0 (camera_module_cache_ram_135__4), .A1 (
          nx36134), .B0 (camera_module_cache_ram_151__4), .B1 (nx36174)) ;
    dffr camera_module_cache_reg_ram_135__4 (.Q (camera_module_cache_ram_135__4)
         , .QB (\$dummy [404]), .D (nx12893), .CLK (clk), .R (rst)) ;
    mux21_ni ix12894 (.Y (nx12893), .A0 (camera_module_cache_ram_135__4), .A1 (
             nx35402), .S0 (nx34612)) ;
    dffr camera_module_cache_reg_ram_151__4 (.Q (camera_module_cache_ram_151__4)
         , .QB (\$dummy [405]), .D (nx12883), .CLK (clk), .R (rst)) ;
    mux21_ni ix12884 (.Y (nx12883), .A0 (camera_module_cache_ram_151__4), .A1 (
             nx35402), .S0 (nx34608)) ;
    aoi22 ix25635 (.Y (nx25634), .A0 (camera_module_cache_ram_183__4), .A1 (
          nx36214), .B0 (camera_module_cache_ram_167__4), .B1 (nx36254)) ;
    dffr camera_module_cache_reg_ram_183__4 (.Q (camera_module_cache_ram_183__4)
         , .QB (\$dummy [406]), .D (nx12863), .CLK (clk), .R (rst)) ;
    mux21_ni ix12864 (.Y (nx12863), .A0 (camera_module_cache_ram_183__4), .A1 (
             nx35402), .S0 (nx34600)) ;
    dffr camera_module_cache_reg_ram_167__4 (.Q (camera_module_cache_ram_167__4)
         , .QB (\$dummy [407]), .D (nx12873), .CLK (clk), .R (rst)) ;
    mux21_ni ix12874 (.Y (nx12873), .A0 (camera_module_cache_ram_167__4), .A1 (
             nx35402), .S0 (nx34604)) ;
    aoi22 ix25645 (.Y (nx25644), .A0 (camera_module_cache_ram_199__4), .A1 (
          nx36294), .B0 (camera_module_cache_ram_215__4), .B1 (nx36334)) ;
    dffr camera_module_cache_reg_ram_199__4 (.Q (camera_module_cache_ram_199__4)
         , .QB (\$dummy [408]), .D (nx12853), .CLK (clk), .R (rst)) ;
    mux21_ni ix12854 (.Y (nx12853), .A0 (camera_module_cache_ram_199__4), .A1 (
             nx35402), .S0 (nx34596)) ;
    dffr camera_module_cache_reg_ram_215__4 (.Q (camera_module_cache_ram_215__4)
         , .QB (\$dummy [409]), .D (nx12843), .CLK (clk), .R (rst)) ;
    mux21_ni ix12844 (.Y (nx12843), .A0 (camera_module_cache_ram_215__4), .A1 (
             nx35402), .S0 (nx34592)) ;
    aoi22 ix25656 (.Y (nx25655), .A0 (camera_module_cache_ram_231__4), .A1 (
          nx36374), .B0 (camera_module_cache_ram_247__4), .B1 (nx36414)) ;
    dffr camera_module_cache_reg_ram_231__4 (.Q (camera_module_cache_ram_231__4)
         , .QB (\$dummy [410]), .D (nx12833), .CLK (clk), .R (rst)) ;
    mux21_ni ix12834 (.Y (nx12833), .A0 (camera_module_cache_ram_231__4), .A1 (
             nx35404), .S0 (nx34588)) ;
    dffr camera_module_cache_reg_ram_247__4 (.Q (camera_module_cache_ram_247__4)
         , .QB (\$dummy [411]), .D (nx12823), .CLK (clk), .R (rst)) ;
    mux21_ni ix12824 (.Y (nx12823), .A0 (camera_module_cache_ram_247__4), .A1 (
             nx35404), .S0 (nx34584)) ;
    nand04 ix15731 (.Y (nx15730), .A0 (nx25667), .A1 (nx25754), .A2 (nx25842), .A3 (
           nx25926)) ;
    oai21 ix25668 (.Y (nx25667), .A0 (nx15720), .A1 (nx15642), .B0 (nx36480)) ;
    nand04 ix15721 (.Y (nx15720), .A0 (nx25671), .A1 (nx25681), .A2 (nx25691), .A3 (
           nx25702)) ;
    aoi22 ix25672 (.Y (nx25671), .A0 (camera_module_cache_ram_8__4), .A1 (
          nx35816), .B0 (camera_module_cache_ram_24__4), .B1 (nx35856)) ;
    dffr camera_module_cache_reg_ram_8__4 (.Q (camera_module_cache_ram_8__4), .QB (
         \$dummy [412]), .D (nx12813), .CLK (clk), .R (rst)) ;
    mux21_ni ix12814 (.Y (nx12813), .A0 (camera_module_cache_ram_8__4), .A1 (
             nx35404), .S0 (nx34574)) ;
    dffr camera_module_cache_reg_ram_24__4 (.Q (camera_module_cache_ram_24__4), 
         .QB (\$dummy [413]), .D (nx12803), .CLK (clk), .R (rst)) ;
    mux21_ni ix12804 (.Y (nx12803), .A0 (camera_module_cache_ram_24__4), .A1 (
             nx35404), .S0 (nx34570)) ;
    aoi22 ix25682 (.Y (nx25681), .A0 (camera_module_cache_ram_40__4), .A1 (
          nx35896), .B0 (camera_module_cache_ram_56__4), .B1 (nx35936)) ;
    dffr camera_module_cache_reg_ram_40__4 (.Q (camera_module_cache_ram_40__4), 
         .QB (\$dummy [414]), .D (nx12793), .CLK (clk), .R (rst)) ;
    mux21_ni ix12794 (.Y (nx12793), .A0 (camera_module_cache_ram_40__4), .A1 (
             nx35404), .S0 (nx34566)) ;
    dffr camera_module_cache_reg_ram_56__4 (.Q (camera_module_cache_ram_56__4), 
         .QB (\$dummy [415]), .D (nx12783), .CLK (clk), .R (rst)) ;
    mux21_ni ix12784 (.Y (nx12783), .A0 (camera_module_cache_ram_56__4), .A1 (
             nx35404), .S0 (nx34562)) ;
    aoi22 ix25692 (.Y (nx25691), .A0 (camera_module_cache_ram_72__4), .A1 (
          nx35976), .B0 (camera_module_cache_ram_88__4), .B1 (nx36016)) ;
    dffr camera_module_cache_reg_ram_72__4 (.Q (camera_module_cache_ram_72__4), 
         .QB (\$dummy [416]), .D (nx12773), .CLK (clk), .R (rst)) ;
    mux21_ni ix12774 (.Y (nx12773), .A0 (camera_module_cache_ram_72__4), .A1 (
             nx35404), .S0 (nx34558)) ;
    dffr camera_module_cache_reg_ram_88__4 (.Q (camera_module_cache_ram_88__4), 
         .QB (\$dummy [417]), .D (nx12763), .CLK (clk), .R (rst)) ;
    mux21_ni ix12764 (.Y (nx12763), .A0 (camera_module_cache_ram_88__4), .A1 (
             nx35406), .S0 (nx34554)) ;
    aoi22 ix25703 (.Y (nx25702), .A0 (camera_module_cache_ram_120__4), .A1 (
          nx36056), .B0 (camera_module_cache_ram_104__4), .B1 (nx36096)) ;
    dffr camera_module_cache_reg_ram_120__4 (.Q (camera_module_cache_ram_120__4)
         , .QB (\$dummy [418]), .D (nx12743), .CLK (clk), .R (rst)) ;
    mux21_ni ix12744 (.Y (nx12743), .A0 (camera_module_cache_ram_120__4), .A1 (
             nx35406), .S0 (nx34546)) ;
    dffr camera_module_cache_reg_ram_104__4 (.Q (camera_module_cache_ram_104__4)
         , .QB (\$dummy [419]), .D (nx12753), .CLK (clk), .R (rst)) ;
    mux21_ni ix12754 (.Y (nx12753), .A0 (camera_module_cache_ram_104__4), .A1 (
             nx35406), .S0 (nx34550)) ;
    nand04 ix15643 (.Y (nx15642), .A0 (nx25711), .A1 (nx25721), .A2 (nx25733), .A3 (
           nx25744)) ;
    aoi22 ix25712 (.Y (nx25711), .A0 (camera_module_cache_ram_136__4), .A1 (
          nx36136), .B0 (camera_module_cache_ram_152__4), .B1 (nx36176)) ;
    dffr camera_module_cache_reg_ram_136__4 (.Q (camera_module_cache_ram_136__4)
         , .QB (\$dummy [420]), .D (nx12733), .CLK (clk), .R (rst)) ;
    mux21_ni ix12734 (.Y (nx12733), .A0 (camera_module_cache_ram_136__4), .A1 (
             nx35406), .S0 (nx34542)) ;
    dffr camera_module_cache_reg_ram_152__4 (.Q (camera_module_cache_ram_152__4)
         , .QB (\$dummy [421]), .D (nx12723), .CLK (clk), .R (rst)) ;
    mux21_ni ix12724 (.Y (nx12723), .A0 (camera_module_cache_ram_152__4), .A1 (
             nx35406), .S0 (nx34538)) ;
    aoi22 ix25722 (.Y (nx25721), .A0 (camera_module_cache_ram_184__4), .A1 (
          nx36216), .B0 (camera_module_cache_ram_168__4), .B1 (nx36256)) ;
    dffr camera_module_cache_reg_ram_184__4 (.Q (camera_module_cache_ram_184__4)
         , .QB (\$dummy [422]), .D (nx12703), .CLK (clk), .R (rst)) ;
    mux21_ni ix12704 (.Y (nx12703), .A0 (camera_module_cache_ram_184__4), .A1 (
             nx35406), .S0 (nx34530)) ;
    dffr camera_module_cache_reg_ram_168__4 (.Q (camera_module_cache_ram_168__4)
         , .QB (\$dummy [423]), .D (nx12713), .CLK (clk), .R (rst)) ;
    mux21_ni ix12714 (.Y (nx12713), .A0 (camera_module_cache_ram_168__4), .A1 (
             nx35406), .S0 (nx34534)) ;
    aoi22 ix25734 (.Y (nx25733), .A0 (camera_module_cache_ram_200__4), .A1 (
          nx36296), .B0 (camera_module_cache_ram_216__4), .B1 (nx36336)) ;
    dffr camera_module_cache_reg_ram_200__4 (.Q (camera_module_cache_ram_200__4)
         , .QB (\$dummy [424]), .D (nx12693), .CLK (clk), .R (rst)) ;
    mux21_ni ix12694 (.Y (nx12693), .A0 (camera_module_cache_ram_200__4), .A1 (
             nx35408), .S0 (nx34526)) ;
    dffr camera_module_cache_reg_ram_216__4 (.Q (camera_module_cache_ram_216__4)
         , .QB (\$dummy [425]), .D (nx12683), .CLK (clk), .R (rst)) ;
    mux21_ni ix12684 (.Y (nx12683), .A0 (camera_module_cache_ram_216__4), .A1 (
             nx35408), .S0 (nx34522)) ;
    aoi22 ix25745 (.Y (nx25744), .A0 (camera_module_cache_ram_232__4), .A1 (
          nx36376), .B0 (camera_module_cache_ram_248__4), .B1 (nx36416)) ;
    dffr camera_module_cache_reg_ram_232__4 (.Q (camera_module_cache_ram_232__4)
         , .QB (\$dummy [426]), .D (nx12673), .CLK (clk), .R (rst)) ;
    mux21_ni ix12674 (.Y (nx12673), .A0 (camera_module_cache_ram_232__4), .A1 (
             nx35408), .S0 (nx34518)) ;
    dffr camera_module_cache_reg_ram_248__4 (.Q (camera_module_cache_ram_248__4)
         , .QB (\$dummy [427]), .D (nx12663), .CLK (clk), .R (rst)) ;
    mux21_ni ix12664 (.Y (nx12663), .A0 (camera_module_cache_ram_248__4), .A1 (
             nx35408), .S0 (nx34514)) ;
    oai21 ix25755 (.Y (nx25754), .A0 (nx15558), .A1 (nx15480), .B0 (nx36484)) ;
    nand04 ix15559 (.Y (nx15558), .A0 (nx25757), .A1 (nx25768), .A2 (nx25778), .A3 (
           nx25787)) ;
    aoi22 ix25758 (.Y (nx25757), .A0 (camera_module_cache_ram_9__4), .A1 (
          nx35816), .B0 (camera_module_cache_ram_25__4), .B1 (nx35856)) ;
    dffr camera_module_cache_reg_ram_9__4 (.Q (camera_module_cache_ram_9__4), .QB (
         \$dummy [428]), .D (nx12653), .CLK (clk), .R (rst)) ;
    mux21_ni ix12654 (.Y (nx12653), .A0 (camera_module_cache_ram_9__4), .A1 (
             nx35408), .S0 (nx34504)) ;
    dffr camera_module_cache_reg_ram_25__4 (.Q (camera_module_cache_ram_25__4), 
         .QB (\$dummy [429]), .D (nx12643), .CLK (clk), .R (rst)) ;
    mux21_ni ix12644 (.Y (nx12643), .A0 (camera_module_cache_ram_25__4), .A1 (
             nx35408), .S0 (nx34500)) ;
    aoi22 ix25769 (.Y (nx25768), .A0 (camera_module_cache_ram_41__4), .A1 (
          nx35896), .B0 (camera_module_cache_ram_57__4), .B1 (nx35936)) ;
    dffr camera_module_cache_reg_ram_41__4 (.Q (camera_module_cache_ram_41__4), 
         .QB (\$dummy [430]), .D (nx12633), .CLK (clk), .R (rst)) ;
    mux21_ni ix12634 (.Y (nx12633), .A0 (camera_module_cache_ram_41__4), .A1 (
             nx35408), .S0 (nx34496)) ;
    dffr camera_module_cache_reg_ram_57__4 (.Q (camera_module_cache_ram_57__4), 
         .QB (\$dummy [431]), .D (nx12623), .CLK (clk), .R (rst)) ;
    mux21_ni ix12624 (.Y (nx12623), .A0 (camera_module_cache_ram_57__4), .A1 (
             nx35410), .S0 (nx34492)) ;
    aoi22 ix25779 (.Y (nx25778), .A0 (camera_module_cache_ram_73__4), .A1 (
          nx35976), .B0 (camera_module_cache_ram_89__4), .B1 (nx36016)) ;
    dffr camera_module_cache_reg_ram_73__4 (.Q (camera_module_cache_ram_73__4), 
         .QB (\$dummy [432]), .D (nx12613), .CLK (clk), .R (rst)) ;
    mux21_ni ix12614 (.Y (nx12613), .A0 (camera_module_cache_ram_73__4), .A1 (
             nx35410), .S0 (nx34488)) ;
    dffr camera_module_cache_reg_ram_89__4 (.Q (camera_module_cache_ram_89__4), 
         .QB (\$dummy [433]), .D (nx12603), .CLK (clk), .R (rst)) ;
    mux21_ni ix12604 (.Y (nx12603), .A0 (camera_module_cache_ram_89__4), .A1 (
             nx35410), .S0 (nx34484)) ;
    aoi22 ix25788 (.Y (nx25787), .A0 (camera_module_cache_ram_121__4), .A1 (
          nx36056), .B0 (camera_module_cache_ram_105__4), .B1 (nx36096)) ;
    dffr camera_module_cache_reg_ram_121__4 (.Q (camera_module_cache_ram_121__4)
         , .QB (\$dummy [434]), .D (nx12583), .CLK (clk), .R (rst)) ;
    mux21_ni ix12584 (.Y (nx12583), .A0 (camera_module_cache_ram_121__4), .A1 (
             nx35410), .S0 (nx34476)) ;
    dffr camera_module_cache_reg_ram_105__4 (.Q (camera_module_cache_ram_105__4)
         , .QB (\$dummy [435]), .D (nx12593), .CLK (clk), .R (rst)) ;
    mux21_ni ix12594 (.Y (nx12593), .A0 (camera_module_cache_ram_105__4), .A1 (
             nx35410), .S0 (nx34480)) ;
    nand04 ix15481 (.Y (nx15480), .A0 (nx25797), .A1 (nx25809), .A2 (nx25821), .A3 (
           nx25831)) ;
    aoi22 ix25798 (.Y (nx25797), .A0 (camera_module_cache_ram_137__4), .A1 (
          nx36136), .B0 (camera_module_cache_ram_153__4), .B1 (nx36176)) ;
    dffr camera_module_cache_reg_ram_137__4 (.Q (camera_module_cache_ram_137__4)
         , .QB (\$dummy [436]), .D (nx12573), .CLK (clk), .R (rst)) ;
    mux21_ni ix12574 (.Y (nx12573), .A0 (camera_module_cache_ram_137__4), .A1 (
             nx35410), .S0 (nx34472)) ;
    dffr camera_module_cache_reg_ram_153__4 (.Q (camera_module_cache_ram_153__4)
         , .QB (\$dummy [437]), .D (nx12563), .CLK (clk), .R (rst)) ;
    mux21_ni ix12564 (.Y (nx12563), .A0 (camera_module_cache_ram_153__4), .A1 (
             nx35410), .S0 (nx34468)) ;
    aoi22 ix25810 (.Y (nx25809), .A0 (camera_module_cache_ram_185__4), .A1 (
          nx36216), .B0 (camera_module_cache_ram_169__4), .B1 (nx36256)) ;
    dffr camera_module_cache_reg_ram_185__4 (.Q (camera_module_cache_ram_185__4)
         , .QB (\$dummy [438]), .D (nx12543), .CLK (clk), .R (rst)) ;
    mux21_ni ix12544 (.Y (nx12543), .A0 (camera_module_cache_ram_185__4), .A1 (
             nx35412), .S0 (nx34460)) ;
    dffr camera_module_cache_reg_ram_169__4 (.Q (camera_module_cache_ram_169__4)
         , .QB (\$dummy [439]), .D (nx12553), .CLK (clk), .R (rst)) ;
    mux21_ni ix12554 (.Y (nx12553), .A0 (camera_module_cache_ram_169__4), .A1 (
             nx35412), .S0 (nx34464)) ;
    aoi22 ix25822 (.Y (nx25821), .A0 (camera_module_cache_ram_201__4), .A1 (
          nx36296), .B0 (camera_module_cache_ram_217__4), .B1 (nx36336)) ;
    dffr camera_module_cache_reg_ram_201__4 (.Q (camera_module_cache_ram_201__4)
         , .QB (\$dummy [440]), .D (nx12533), .CLK (clk), .R (rst)) ;
    mux21_ni ix12534 (.Y (nx12533), .A0 (camera_module_cache_ram_201__4), .A1 (
             nx35412), .S0 (nx34456)) ;
    dffr camera_module_cache_reg_ram_217__4 (.Q (camera_module_cache_ram_217__4)
         , .QB (\$dummy [441]), .D (nx12523), .CLK (clk), .R (rst)) ;
    mux21_ni ix12524 (.Y (nx12523), .A0 (camera_module_cache_ram_217__4), .A1 (
             nx35412), .S0 (nx34452)) ;
    aoi22 ix25832 (.Y (nx25831), .A0 (camera_module_cache_ram_233__4), .A1 (
          nx36376), .B0 (camera_module_cache_ram_249__4), .B1 (nx36416)) ;
    dffr camera_module_cache_reg_ram_233__4 (.Q (camera_module_cache_ram_233__4)
         , .QB (\$dummy [442]), .D (nx12513), .CLK (clk), .R (rst)) ;
    mux21_ni ix12514 (.Y (nx12513), .A0 (camera_module_cache_ram_233__4), .A1 (
             nx35412), .S0 (nx34448)) ;
    dffr camera_module_cache_reg_ram_249__4 (.Q (camera_module_cache_ram_249__4)
         , .QB (\$dummy [443]), .D (nx12503), .CLK (clk), .R (rst)) ;
    mux21_ni ix12504 (.Y (nx12503), .A0 (camera_module_cache_ram_249__4), .A1 (
             nx35412), .S0 (nx34444)) ;
    oai21 ix25843 (.Y (nx25842), .A0 (nx15394), .A1 (nx15316), .B0 (nx36488)) ;
    nand04 ix15395 (.Y (nx15394), .A0 (nx25845), .A1 (nx25855), .A2 (nx25864), .A3 (
           nx25872)) ;
    aoi22 ix25846 (.Y (nx25845), .A0 (camera_module_cache_ram_10__4), .A1 (
          nx35816), .B0 (camera_module_cache_ram_26__4), .B1 (nx35856)) ;
    dffr camera_module_cache_reg_ram_10__4 (.Q (camera_module_cache_ram_10__4), 
         .QB (\$dummy [444]), .D (nx12493), .CLK (clk), .R (rst)) ;
    mux21_ni ix12494 (.Y (nx12493), .A0 (camera_module_cache_ram_10__4), .A1 (
             nx35412), .S0 (nx34434)) ;
    dffr camera_module_cache_reg_ram_26__4 (.Q (camera_module_cache_ram_26__4), 
         .QB (\$dummy [445]), .D (nx12483), .CLK (clk), .R (rst)) ;
    mux21_ni ix12484 (.Y (nx12483), .A0 (camera_module_cache_ram_26__4), .A1 (
             nx35414), .S0 (nx34430)) ;
    aoi22 ix25856 (.Y (nx25855), .A0 (camera_module_cache_ram_42__4), .A1 (
          nx35896), .B0 (camera_module_cache_ram_58__4), .B1 (nx35936)) ;
    dffr camera_module_cache_reg_ram_42__4 (.Q (camera_module_cache_ram_42__4), 
         .QB (\$dummy [446]), .D (nx12473), .CLK (clk), .R (rst)) ;
    mux21_ni ix12474 (.Y (nx12473), .A0 (camera_module_cache_ram_42__4), .A1 (
             nx35414), .S0 (nx34426)) ;
    dffr camera_module_cache_reg_ram_58__4 (.Q (camera_module_cache_ram_58__4), 
         .QB (\$dummy [447]), .D (nx12463), .CLK (clk), .R (rst)) ;
    mux21_ni ix12464 (.Y (nx12463), .A0 (camera_module_cache_ram_58__4), .A1 (
             nx35414), .S0 (nx34422)) ;
    aoi22 ix25865 (.Y (nx25864), .A0 (camera_module_cache_ram_74__4), .A1 (
          nx35976), .B0 (camera_module_cache_ram_90__4), .B1 (nx36016)) ;
    dffr camera_module_cache_reg_ram_74__4 (.Q (camera_module_cache_ram_74__4), 
         .QB (\$dummy [448]), .D (nx12453), .CLK (clk), .R (rst)) ;
    mux21_ni ix12454 (.Y (nx12453), .A0 (camera_module_cache_ram_74__4), .A1 (
             nx35414), .S0 (nx34418)) ;
    dffr camera_module_cache_reg_ram_90__4 (.Q (camera_module_cache_ram_90__4), 
         .QB (\$dummy [449]), .D (nx12443), .CLK (clk), .R (rst)) ;
    mux21_ni ix12444 (.Y (nx12443), .A0 (camera_module_cache_ram_90__4), .A1 (
             nx35414), .S0 (nx34414)) ;
    aoi22 ix25874 (.Y (nx25872), .A0 (camera_module_cache_ram_122__4), .A1 (
          nx36056), .B0 (camera_module_cache_ram_106__4), .B1 (nx36096)) ;
    dffr camera_module_cache_reg_ram_122__4 (.Q (camera_module_cache_ram_122__4)
         , .QB (\$dummy [450]), .D (nx12423), .CLK (clk), .R (rst)) ;
    mux21_ni ix12424 (.Y (nx12423), .A0 (camera_module_cache_ram_122__4), .A1 (
             nx35414), .S0 (nx34406)) ;
    dffr camera_module_cache_reg_ram_106__4 (.Q (camera_module_cache_ram_106__4)
         , .QB (\$dummy [451]), .D (nx12433), .CLK (clk), .R (rst)) ;
    mux21_ni ix12434 (.Y (nx12433), .A0 (camera_module_cache_ram_106__4), .A1 (
             nx35414), .S0 (nx34410)) ;
    nand04 ix15317 (.Y (nx15316), .A0 (nx25885), .A1 (nx25895), .A2 (nx25905), .A3 (
           nx25916)) ;
    aoi22 ix25886 (.Y (nx25885), .A0 (camera_module_cache_ram_138__4), .A1 (
          nx36136), .B0 (camera_module_cache_ram_154__4), .B1 (nx36176)) ;
    dffr camera_module_cache_reg_ram_138__4 (.Q (camera_module_cache_ram_138__4)
         , .QB (\$dummy [452]), .D (nx12413), .CLK (clk), .R (rst)) ;
    mux21_ni ix12414 (.Y (nx12413), .A0 (camera_module_cache_ram_138__4), .A1 (
             nx35416), .S0 (nx34402)) ;
    dffr camera_module_cache_reg_ram_154__4 (.Q (camera_module_cache_ram_154__4)
         , .QB (\$dummy [453]), .D (nx12403), .CLK (clk), .R (rst)) ;
    mux21_ni ix12404 (.Y (nx12403), .A0 (camera_module_cache_ram_154__4), .A1 (
             nx35416), .S0 (nx34398)) ;
    aoi22 ix25896 (.Y (nx25895), .A0 (camera_module_cache_ram_186__4), .A1 (
          nx36216), .B0 (camera_module_cache_ram_170__4), .B1 (nx36256)) ;
    dffr camera_module_cache_reg_ram_186__4 (.Q (camera_module_cache_ram_186__4)
         , .QB (\$dummy [454]), .D (nx12383), .CLK (clk), .R (rst)) ;
    mux21_ni ix12384 (.Y (nx12383), .A0 (camera_module_cache_ram_186__4), .A1 (
             nx35416), .S0 (nx34390)) ;
    dffr camera_module_cache_reg_ram_170__4 (.Q (camera_module_cache_ram_170__4)
         , .QB (\$dummy [455]), .D (nx12393), .CLK (clk), .R (rst)) ;
    mux21_ni ix12394 (.Y (nx12393), .A0 (camera_module_cache_ram_170__4), .A1 (
             nx35416), .S0 (nx34394)) ;
    aoi22 ix25906 (.Y (nx25905), .A0 (camera_module_cache_ram_202__4), .A1 (
          nx36296), .B0 (camera_module_cache_ram_218__4), .B1 (nx36336)) ;
    dffr camera_module_cache_reg_ram_202__4 (.Q (camera_module_cache_ram_202__4)
         , .QB (\$dummy [456]), .D (nx12373), .CLK (clk), .R (rst)) ;
    mux21_ni ix12374 (.Y (nx12373), .A0 (camera_module_cache_ram_202__4), .A1 (
             nx35416), .S0 (nx34386)) ;
    dffr camera_module_cache_reg_ram_218__4 (.Q (camera_module_cache_ram_218__4)
         , .QB (\$dummy [457]), .D (nx12363), .CLK (clk), .R (rst)) ;
    mux21_ni ix12364 (.Y (nx12363), .A0 (camera_module_cache_ram_218__4), .A1 (
             nx35416), .S0 (nx34382)) ;
    aoi22 ix25917 (.Y (nx25916), .A0 (camera_module_cache_ram_234__4), .A1 (
          nx36376), .B0 (camera_module_cache_ram_250__4), .B1 (nx36416)) ;
    dffr camera_module_cache_reg_ram_234__4 (.Q (camera_module_cache_ram_234__4)
         , .QB (\$dummy [458]), .D (nx12353), .CLK (clk), .R (rst)) ;
    mux21_ni ix12354 (.Y (nx12353), .A0 (camera_module_cache_ram_234__4), .A1 (
             nx35416), .S0 (nx34378)) ;
    dffr camera_module_cache_reg_ram_250__4 (.Q (camera_module_cache_ram_250__4)
         , .QB (\$dummy [459]), .D (nx12343), .CLK (clk), .R (rst)) ;
    mux21_ni ix12344 (.Y (nx12343), .A0 (camera_module_cache_ram_250__4), .A1 (
             nx35418), .S0 (nx34374)) ;
    oai21 ix25927 (.Y (nx25926), .A0 (nx15232), .A1 (nx15154), .B0 (nx36492)) ;
    nand04 ix15233 (.Y (nx15232), .A0 (nx25929), .A1 (nx25938), .A2 (nx25946), .A3 (
           nx25959)) ;
    aoi22 ix25930 (.Y (nx25929), .A0 (camera_module_cache_ram_11__4), .A1 (
          nx35816), .B0 (camera_module_cache_ram_27__4), .B1 (nx35856)) ;
    dffr camera_module_cache_reg_ram_11__4 (.Q (camera_module_cache_ram_11__4), 
         .QB (\$dummy [460]), .D (nx12333), .CLK (clk), .R (rst)) ;
    mux21_ni ix12334 (.Y (nx12333), .A0 (camera_module_cache_ram_11__4), .A1 (
             nx35418), .S0 (nx34364)) ;
    dffr camera_module_cache_reg_ram_27__4 (.Q (camera_module_cache_ram_27__4), 
         .QB (\$dummy [461]), .D (nx12323), .CLK (clk), .R (rst)) ;
    mux21_ni ix12324 (.Y (nx12323), .A0 (camera_module_cache_ram_27__4), .A1 (
             nx35418), .S0 (nx34360)) ;
    aoi22 ix25939 (.Y (nx25938), .A0 (camera_module_cache_ram_43__4), .A1 (
          nx35896), .B0 (camera_module_cache_ram_59__4), .B1 (nx35936)) ;
    dffr camera_module_cache_reg_ram_43__4 (.Q (camera_module_cache_ram_43__4), 
         .QB (\$dummy [462]), .D (nx12313), .CLK (clk), .R (rst)) ;
    mux21_ni ix12314 (.Y (nx12313), .A0 (camera_module_cache_ram_43__4), .A1 (
             nx35418), .S0 (nx34356)) ;
    dffr camera_module_cache_reg_ram_59__4 (.Q (camera_module_cache_ram_59__4), 
         .QB (\$dummy [463]), .D (nx12303), .CLK (clk), .R (rst)) ;
    mux21_ni ix12304 (.Y (nx12303), .A0 (camera_module_cache_ram_59__4), .A1 (
             nx35418), .S0 (nx34352)) ;
    aoi22 ix25948 (.Y (nx25946), .A0 (camera_module_cache_ram_75__4), .A1 (
          nx35976), .B0 (camera_module_cache_ram_91__4), .B1 (nx36016)) ;
    dffr camera_module_cache_reg_ram_75__4 (.Q (camera_module_cache_ram_75__4), 
         .QB (\$dummy [464]), .D (nx12293), .CLK (clk), .R (rst)) ;
    mux21_ni ix12294 (.Y (nx12293), .A0 (camera_module_cache_ram_75__4), .A1 (
             nx35418), .S0 (nx34348)) ;
    dffr camera_module_cache_reg_ram_91__4 (.Q (camera_module_cache_ram_91__4), 
         .QB (\$dummy [465]), .D (nx12283), .CLK (clk), .R (rst)) ;
    mux21_ni ix12284 (.Y (nx12283), .A0 (camera_module_cache_ram_91__4), .A1 (
             nx35418), .S0 (nx34344)) ;
    aoi22 ix25960 (.Y (nx25959), .A0 (camera_module_cache_ram_123__4), .A1 (
          nx36056), .B0 (camera_module_cache_ram_107__4), .B1 (nx36096)) ;
    dffr camera_module_cache_reg_ram_123__4 (.Q (camera_module_cache_ram_123__4)
         , .QB (\$dummy [466]), .D (nx12263), .CLK (clk), .R (rst)) ;
    mux21_ni ix12264 (.Y (nx12263), .A0 (camera_module_cache_ram_123__4), .A1 (
             nx35420), .S0 (nx34336)) ;
    dffr camera_module_cache_reg_ram_107__4 (.Q (camera_module_cache_ram_107__4)
         , .QB (\$dummy [467]), .D (nx12273), .CLK (clk), .R (rst)) ;
    mux21_ni ix12274 (.Y (nx12273), .A0 (camera_module_cache_ram_107__4), .A1 (
             nx35420), .S0 (nx34340)) ;
    nand04 ix15155 (.Y (nx15154), .A0 (nx25969), .A1 (nx25979), .A2 (nx25990), .A3 (
           nx26000)) ;
    aoi22 ix25970 (.Y (nx25969), .A0 (camera_module_cache_ram_139__4), .A1 (
          nx36136), .B0 (camera_module_cache_ram_155__4), .B1 (nx36176)) ;
    dffr camera_module_cache_reg_ram_139__4 (.Q (camera_module_cache_ram_139__4)
         , .QB (\$dummy [468]), .D (nx12253), .CLK (clk), .R (rst)) ;
    mux21_ni ix12254 (.Y (nx12253), .A0 (camera_module_cache_ram_139__4), .A1 (
             nx35420), .S0 (nx34332)) ;
    dffr camera_module_cache_reg_ram_155__4 (.Q (camera_module_cache_ram_155__4)
         , .QB (\$dummy [469]), .D (nx12243), .CLK (clk), .R (rst)) ;
    mux21_ni ix12244 (.Y (nx12243), .A0 (camera_module_cache_ram_155__4), .A1 (
             nx35420), .S0 (nx34328)) ;
    aoi22 ix25980 (.Y (nx25979), .A0 (camera_module_cache_ram_187__4), .A1 (
          nx36216), .B0 (camera_module_cache_ram_171__4), .B1 (nx36256)) ;
    dffr camera_module_cache_reg_ram_187__4 (.Q (camera_module_cache_ram_187__4)
         , .QB (\$dummy [470]), .D (nx12223), .CLK (clk), .R (rst)) ;
    mux21_ni ix12224 (.Y (nx12223), .A0 (camera_module_cache_ram_187__4), .A1 (
             nx35420), .S0 (nx34320)) ;
    dffr camera_module_cache_reg_ram_171__4 (.Q (camera_module_cache_ram_171__4)
         , .QB (\$dummy [471]), .D (nx12233), .CLK (clk), .R (rst)) ;
    mux21_ni ix12234 (.Y (nx12233), .A0 (camera_module_cache_ram_171__4), .A1 (
             nx35420), .S0 (nx34324)) ;
    aoi22 ix25991 (.Y (nx25990), .A0 (camera_module_cache_ram_203__4), .A1 (
          nx36296), .B0 (camera_module_cache_ram_219__4), .B1 (nx36336)) ;
    dffr camera_module_cache_reg_ram_203__4 (.Q (camera_module_cache_ram_203__4)
         , .QB (\$dummy [472]), .D (nx12213), .CLK (clk), .R (rst)) ;
    mux21_ni ix12214 (.Y (nx12213), .A0 (camera_module_cache_ram_203__4), .A1 (
             nx35420), .S0 (nx34316)) ;
    dffr camera_module_cache_reg_ram_219__4 (.Q (camera_module_cache_ram_219__4)
         , .QB (\$dummy [473]), .D (nx12203), .CLK (clk), .R (rst)) ;
    mux21_ni ix12204 (.Y (nx12203), .A0 (camera_module_cache_ram_219__4), .A1 (
             nx35422), .S0 (nx34312)) ;
    aoi22 ix26001 (.Y (nx26000), .A0 (camera_module_cache_ram_235__4), .A1 (
          nx36376), .B0 (camera_module_cache_ram_251__4), .B1 (nx36416)) ;
    dffr camera_module_cache_reg_ram_235__4 (.Q (camera_module_cache_ram_235__4)
         , .QB (\$dummy [474]), .D (nx12193), .CLK (clk), .R (rst)) ;
    mux21_ni ix12194 (.Y (nx12193), .A0 (camera_module_cache_ram_235__4), .A1 (
             nx35422), .S0 (nx34308)) ;
    dffr camera_module_cache_reg_ram_251__4 (.Q (camera_module_cache_ram_251__4)
         , .QB (\$dummy [475]), .D (nx12183), .CLK (clk), .R (rst)) ;
    mux21_ni ix12184 (.Y (nx12183), .A0 (camera_module_cache_ram_251__4), .A1 (
             nx35422), .S0 (nx34304)) ;
    nand04 ix15077 (.Y (nx15076), .A0 (nx26009), .A1 (nx26094), .A2 (nx26185), .A3 (
           nx26272)) ;
    oai21 ix26010 (.Y (nx26009), .A0 (nx15066), .A1 (nx14988), .B0 (nx36506)) ;
    nand04 ix15067 (.Y (nx15066), .A0 (nx26013), .A1 (nx26023), .A2 (nx26034), .A3 (
           nx26045)) ;
    aoi22 ix26014 (.Y (nx26013), .A0 (camera_module_cache_ram_12__4), .A1 (
          nx35816), .B0 (camera_module_cache_ram_28__4), .B1 (nx35856)) ;
    dffr camera_module_cache_reg_ram_12__4 (.Q (camera_module_cache_ram_12__4), 
         .QB (\$dummy [476]), .D (nx12173), .CLK (clk), .R (rst)) ;
    mux21_ni ix12174 (.Y (nx12173), .A0 (nx35422), .A1 (
             camera_module_cache_ram_12__4), .S0 (nx36496)) ;
    dffr camera_module_cache_reg_ram_28__4 (.Q (camera_module_cache_ram_28__4), 
         .QB (\$dummy [477]), .D (nx12163), .CLK (clk), .R (rst)) ;
    mux21_ni ix12164 (.Y (nx12163), .A0 (nx35422), .A1 (
             camera_module_cache_ram_28__4), .S0 (nx36510)) ;
    aoi22 ix26024 (.Y (nx26023), .A0 (camera_module_cache_ram_44__4), .A1 (
          nx35896), .B0 (camera_module_cache_ram_60__4), .B1 (nx35936)) ;
    dffr camera_module_cache_reg_ram_44__4 (.Q (camera_module_cache_ram_44__4), 
         .QB (\$dummy [478]), .D (nx12153), .CLK (clk), .R (rst)) ;
    mux21_ni ix12154 (.Y (nx12153), .A0 (nx35422), .A1 (
             camera_module_cache_ram_44__4), .S0 (nx36514)) ;
    dffr camera_module_cache_reg_ram_60__4 (.Q (camera_module_cache_ram_60__4), 
         .QB (\$dummy [479]), .D (nx12143), .CLK (clk), .R (rst)) ;
    mux21_ni ix12144 (.Y (nx12143), .A0 (nx35422), .A1 (
             camera_module_cache_ram_60__4), .S0 (nx36518)) ;
    aoi22 ix26035 (.Y (nx26034), .A0 (camera_module_cache_ram_76__4), .A1 (
          nx35976), .B0 (camera_module_cache_ram_92__4), .B1 (nx36016)) ;
    dffr camera_module_cache_reg_ram_76__4 (.Q (camera_module_cache_ram_76__4), 
         .QB (\$dummy [480]), .D (nx12133), .CLK (clk), .R (rst)) ;
    mux21_ni ix12134 (.Y (nx12133), .A0 (nx35424), .A1 (
             camera_module_cache_ram_76__4), .S0 (nx36522)) ;
    dffr camera_module_cache_reg_ram_92__4 (.Q (camera_module_cache_ram_92__4), 
         .QB (\$dummy [481]), .D (nx12123), .CLK (clk), .R (rst)) ;
    mux21_ni ix12124 (.Y (nx12123), .A0 (nx35424), .A1 (
             camera_module_cache_ram_92__4), .S0 (nx36526)) ;
    aoi22 ix26046 (.Y (nx26045), .A0 (camera_module_cache_ram_124__4), .A1 (
          nx36056), .B0 (camera_module_cache_ram_108__4), .B1 (nx36096)) ;
    dffr camera_module_cache_reg_ram_124__4 (.Q (camera_module_cache_ram_124__4)
         , .QB (\$dummy [482]), .D (nx12103), .CLK (clk), .R (rst)) ;
    mux21_ni ix12104 (.Y (nx12103), .A0 (nx35424), .A1 (
             camera_module_cache_ram_124__4), .S0 (nx36530)) ;
    dffr camera_module_cache_reg_ram_108__4 (.Q (camera_module_cache_ram_108__4)
         , .QB (\$dummy [483]), .D (nx12113), .CLK (clk), .R (rst)) ;
    mux21_ni ix12114 (.Y (nx12113), .A0 (nx35424), .A1 (
             camera_module_cache_ram_108__4), .S0 (nx36534)) ;
    nand04 ix14989 (.Y (nx14988), .A0 (nx26055), .A1 (nx26067), .A2 (nx26077), .A3 (
           nx26086)) ;
    aoi22 ix26056 (.Y (nx26055), .A0 (camera_module_cache_ram_140__4), .A1 (
          nx36136), .B0 (camera_module_cache_ram_156__4), .B1 (nx36176)) ;
    dffr camera_module_cache_reg_ram_140__4 (.Q (camera_module_cache_ram_140__4)
         , .QB (\$dummy [484]), .D (nx12093), .CLK (clk), .R (rst)) ;
    mux21_ni ix12094 (.Y (nx12093), .A0 (nx35424), .A1 (
             camera_module_cache_ram_140__4), .S0 (nx36538)) ;
    dffr camera_module_cache_reg_ram_156__4 (.Q (camera_module_cache_ram_156__4)
         , .QB (\$dummy [485]), .D (nx12083), .CLK (clk), .R (rst)) ;
    mux21_ni ix12084 (.Y (nx12083), .A0 (nx35424), .A1 (
             camera_module_cache_ram_156__4), .S0 (nx36542)) ;
    aoi22 ix26068 (.Y (nx26067), .A0 (camera_module_cache_ram_188__4), .A1 (
          nx36216), .B0 (camera_module_cache_ram_172__4), .B1 (nx36256)) ;
    dffr camera_module_cache_reg_ram_188__4 (.Q (camera_module_cache_ram_188__4)
         , .QB (\$dummy [486]), .D (nx12063), .CLK (clk), .R (rst)) ;
    mux21_ni ix12064 (.Y (nx12063), .A0 (nx35424), .A1 (
             camera_module_cache_ram_188__4), .S0 (nx36546)) ;
    dffr camera_module_cache_reg_ram_172__4 (.Q (camera_module_cache_ram_172__4)
         , .QB (\$dummy [487]), .D (nx12073), .CLK (clk), .R (rst)) ;
    mux21_ni ix12074 (.Y (nx12073), .A0 (nx35426), .A1 (
             camera_module_cache_ram_172__4), .S0 (nx36550)) ;
    aoi22 ix26078 (.Y (nx26077), .A0 (camera_module_cache_ram_204__4), .A1 (
          nx36296), .B0 (camera_module_cache_ram_220__4), .B1 (nx36336)) ;
    dffr camera_module_cache_reg_ram_204__4 (.Q (camera_module_cache_ram_204__4)
         , .QB (\$dummy [488]), .D (nx12053), .CLK (clk), .R (rst)) ;
    mux21_ni ix12054 (.Y (nx12053), .A0 (nx35426), .A1 (
             camera_module_cache_ram_204__4), .S0 (nx36554)) ;
    dffr camera_module_cache_reg_ram_220__4 (.Q (camera_module_cache_ram_220__4)
         , .QB (\$dummy [489]), .D (nx12043), .CLK (clk), .R (rst)) ;
    mux21_ni ix12044 (.Y (nx12043), .A0 (nx35426), .A1 (
             camera_module_cache_ram_220__4), .S0 (nx36558)) ;
    aoi22 ix26087 (.Y (nx26086), .A0 (camera_module_cache_ram_236__4), .A1 (
          nx36376), .B0 (camera_module_cache_ram_252__4), .B1 (nx36416)) ;
    dffr camera_module_cache_reg_ram_236__4 (.Q (camera_module_cache_ram_236__4)
         , .QB (\$dummy [490]), .D (nx12033), .CLK (clk), .R (rst)) ;
    mux21_ni ix12034 (.Y (nx12033), .A0 (nx35426), .A1 (
             camera_module_cache_ram_236__4), .S0 (nx36562)) ;
    dffr camera_module_cache_reg_ram_252__4 (.Q (camera_module_cache_ram_252__4)
         , .QB (\$dummy [491]), .D (nx12023), .CLK (clk), .R (rst)) ;
    mux21_ni ix12024 (.Y (nx12023), .A0 (nx35426), .A1 (
             camera_module_cache_ram_252__4), .S0 (nx36566)) ;
    oai21 ix26096 (.Y (nx26094), .A0 (nx14904), .A1 (nx14826), .B0 (nx36580)) ;
    nand04 ix14905 (.Y (nx14904), .A0 (nx26099), .A1 (nx26111), .A2 (nx26122), .A3 (
           nx26131)) ;
    aoi22 ix26100 (.Y (nx26099), .A0 (camera_module_cache_ram_13__4), .A1 (
          nx35816), .B0 (camera_module_cache_ram_29__4), .B1 (nx35856)) ;
    dffr camera_module_cache_reg_ram_13__4 (.Q (camera_module_cache_ram_13__4), 
         .QB (\$dummy [492]), .D (nx12013), .CLK (clk), .R (rst)) ;
    mux21_ni ix12014 (.Y (nx12013), .A0 (nx35426), .A1 (
             camera_module_cache_ram_13__4), .S0 (nx36570)) ;
    dffr camera_module_cache_reg_ram_29__4 (.Q (camera_module_cache_ram_29__4), 
         .QB (\$dummy [493]), .D (nx12003), .CLK (clk), .R (rst)) ;
    mux21_ni ix12004 (.Y (nx12003), .A0 (nx35426), .A1 (
             camera_module_cache_ram_29__4), .S0 (nx36584)) ;
    aoi22 ix26112 (.Y (nx26111), .A0 (camera_module_cache_ram_45__4), .A1 (
          nx35896), .B0 (camera_module_cache_ram_61__4), .B1 (nx35936)) ;
    dffr camera_module_cache_reg_ram_45__4 (.Q (camera_module_cache_ram_45__4), 
         .QB (\$dummy [494]), .D (nx11993), .CLK (clk), .R (rst)) ;
    mux21_ni ix11994 (.Y (nx11993), .A0 (nx35428), .A1 (
             camera_module_cache_ram_45__4), .S0 (nx36588)) ;
    dffr camera_module_cache_reg_ram_61__4 (.Q (camera_module_cache_ram_61__4), 
         .QB (\$dummy [495]), .D (nx11983), .CLK (clk), .R (rst)) ;
    mux21_ni ix11984 (.Y (nx11983), .A0 (nx35428), .A1 (
             camera_module_cache_ram_61__4), .S0 (nx36592)) ;
    aoi22 ix26123 (.Y (nx26122), .A0 (camera_module_cache_ram_77__4), .A1 (
          nx35976), .B0 (camera_module_cache_ram_93__4), .B1 (nx36016)) ;
    dffr camera_module_cache_reg_ram_77__4 (.Q (camera_module_cache_ram_77__4), 
         .QB (\$dummy [496]), .D (nx11973), .CLK (clk), .R (rst)) ;
    mux21_ni ix11974 (.Y (nx11973), .A0 (nx35428), .A1 (
             camera_module_cache_ram_77__4), .S0 (nx36596)) ;
    dffr camera_module_cache_reg_ram_93__4 (.Q (camera_module_cache_ram_93__4), 
         .QB (\$dummy [497]), .D (nx11963), .CLK (clk), .R (rst)) ;
    mux21_ni ix11964 (.Y (nx11963), .A0 (nx35428), .A1 (
             camera_module_cache_ram_93__4), .S0 (nx36600)) ;
    aoi22 ix26132 (.Y (nx26131), .A0 (camera_module_cache_ram_125__4), .A1 (
          nx36056), .B0 (camera_module_cache_ram_109__4), .B1 (nx36096)) ;
    dffr camera_module_cache_reg_ram_125__4 (.Q (camera_module_cache_ram_125__4)
         , .QB (\$dummy [498]), .D (nx11943), .CLK (clk), .R (rst)) ;
    mux21_ni ix11944 (.Y (nx11943), .A0 (nx35428), .A1 (
             camera_module_cache_ram_125__4), .S0 (nx36604)) ;
    dffr camera_module_cache_reg_ram_109__4 (.Q (camera_module_cache_ram_109__4)
         , .QB (\$dummy [499]), .D (nx11953), .CLK (clk), .R (rst)) ;
    mux21_ni ix11954 (.Y (nx11953), .A0 (nx35428), .A1 (
             camera_module_cache_ram_109__4), .S0 (nx36608)) ;
    nand04 ix14827 (.Y (nx14826), .A0 (nx26143), .A1 (nx26152), .A2 (nx26162), .A3 (
           nx26173)) ;
    aoi22 ix26144 (.Y (nx26143), .A0 (camera_module_cache_ram_141__4), .A1 (
          nx36136), .B0 (camera_module_cache_ram_157__4), .B1 (nx36176)) ;
    dffr camera_module_cache_reg_ram_141__4 (.Q (camera_module_cache_ram_141__4)
         , .QB (\$dummy [500]), .D (nx11933), .CLK (clk), .R (rst)) ;
    mux21_ni ix11934 (.Y (nx11933), .A0 (nx35428), .A1 (
             camera_module_cache_ram_141__4), .S0 (nx36612)) ;
    dffr camera_module_cache_reg_ram_157__4 (.Q (camera_module_cache_ram_157__4)
         , .QB (\$dummy [501]), .D (nx11923), .CLK (clk), .R (rst)) ;
    mux21_ni ix11924 (.Y (nx11923), .A0 (nx35430), .A1 (
             camera_module_cache_ram_157__4), .S0 (nx36616)) ;
    aoi22 ix26153 (.Y (nx26152), .A0 (camera_module_cache_ram_189__4), .A1 (
          nx36216), .B0 (camera_module_cache_ram_173__4), .B1 (nx36256)) ;
    dffr camera_module_cache_reg_ram_189__4 (.Q (camera_module_cache_ram_189__4)
         , .QB (\$dummy [502]), .D (nx11903), .CLK (clk), .R (rst)) ;
    mux21_ni ix11904 (.Y (nx11903), .A0 (nx35430), .A1 (
             camera_module_cache_ram_189__4), .S0 (nx36620)) ;
    dffr camera_module_cache_reg_ram_173__4 (.Q (camera_module_cache_ram_173__4)
         , .QB (\$dummy [503]), .D (nx11913), .CLK (clk), .R (rst)) ;
    mux21_ni ix11914 (.Y (nx11913), .A0 (nx35430), .A1 (
             camera_module_cache_ram_173__4), .S0 (nx36624)) ;
    aoi22 ix26163 (.Y (nx26162), .A0 (camera_module_cache_ram_205__4), .A1 (
          nx36296), .B0 (camera_module_cache_ram_221__4), .B1 (nx36336)) ;
    dffr camera_module_cache_reg_ram_205__4 (.Q (camera_module_cache_ram_205__4)
         , .QB (\$dummy [504]), .D (nx11893), .CLK (clk), .R (rst)) ;
    mux21_ni ix11894 (.Y (nx11893), .A0 (nx35430), .A1 (
             camera_module_cache_ram_205__4), .S0 (nx36628)) ;
    dffr camera_module_cache_reg_ram_221__4 (.Q (camera_module_cache_ram_221__4)
         , .QB (\$dummy [505]), .D (nx11883), .CLK (clk), .R (rst)) ;
    mux21_ni ix11884 (.Y (nx11883), .A0 (nx35430), .A1 (
             camera_module_cache_ram_221__4), .S0 (nx36632)) ;
    aoi22 ix26174 (.Y (nx26173), .A0 (camera_module_cache_ram_237__4), .A1 (
          nx36376), .B0 (camera_module_cache_ram_253__4), .B1 (nx36416)) ;
    dffr camera_module_cache_reg_ram_237__4 (.Q (camera_module_cache_ram_237__4)
         , .QB (\$dummy [506]), .D (nx11873), .CLK (clk), .R (rst)) ;
    mux21_ni ix11874 (.Y (nx11873), .A0 (nx35430), .A1 (
             camera_module_cache_ram_237__4), .S0 (nx36636)) ;
    dffr camera_module_cache_reg_ram_253__4 (.Q (camera_module_cache_ram_253__4)
         , .QB (\$dummy [507]), .D (nx11863), .CLK (clk), .R (rst)) ;
    mux21_ni ix11864 (.Y (nx11863), .A0 (nx35430), .A1 (
             camera_module_cache_ram_253__4), .S0 (nx36640)) ;
    oai21 ix26186 (.Y (nx26185), .A0 (nx14740), .A1 (nx14662), .B0 (nx36654)) ;
    nand04 ix14741 (.Y (nx14740), .A0 (nx26189), .A1 (nx26199), .A2 (nx26209), .A3 (
           nx26220)) ;
    aoi22 ix26190 (.Y (nx26189), .A0 (camera_module_cache_ram_14__4), .A1 (
          nx35816), .B0 (camera_module_cache_ram_30__4), .B1 (nx35856)) ;
    dffr camera_module_cache_reg_ram_14__4 (.Q (camera_module_cache_ram_14__4), 
         .QB (\$dummy [508]), .D (nx11853), .CLK (clk), .R (rst)) ;
    mux21_ni ix11854 (.Y (nx11853), .A0 (nx35432), .A1 (
             camera_module_cache_ram_14__4), .S0 (nx36644)) ;
    dffr camera_module_cache_reg_ram_30__4 (.Q (camera_module_cache_ram_30__4), 
         .QB (\$dummy [509]), .D (nx11843), .CLK (clk), .R (rst)) ;
    mux21_ni ix11844 (.Y (nx11843), .A0 (nx35432), .A1 (
             camera_module_cache_ram_30__4), .S0 (nx36658)) ;
    aoi22 ix26200 (.Y (nx26199), .A0 (camera_module_cache_ram_46__4), .A1 (
          nx35896), .B0 (camera_module_cache_ram_62__4), .B1 (nx35936)) ;
    dffr camera_module_cache_reg_ram_46__4 (.Q (camera_module_cache_ram_46__4), 
         .QB (\$dummy [510]), .D (nx11833), .CLK (clk), .R (rst)) ;
    mux21_ni ix11834 (.Y (nx11833), .A0 (nx35432), .A1 (
             camera_module_cache_ram_46__4), .S0 (nx36662)) ;
    dffr camera_module_cache_reg_ram_62__4 (.Q (camera_module_cache_ram_62__4), 
         .QB (\$dummy [511]), .D (nx11823), .CLK (clk), .R (rst)) ;
    mux21_ni ix11824 (.Y (nx11823), .A0 (nx35432), .A1 (
             camera_module_cache_ram_62__4), .S0 (nx36666)) ;
    aoi22 ix26210 (.Y (nx26209), .A0 (camera_module_cache_ram_78__4), .A1 (
          nx35976), .B0 (camera_module_cache_ram_94__4), .B1 (nx36016)) ;
    dffr camera_module_cache_reg_ram_78__4 (.Q (camera_module_cache_ram_78__4), 
         .QB (\$dummy [512]), .D (nx11813), .CLK (clk), .R (rst)) ;
    mux21_ni ix11814 (.Y (nx11813), .A0 (nx35432), .A1 (
             camera_module_cache_ram_78__4), .S0 (nx36670)) ;
    dffr camera_module_cache_reg_ram_94__4 (.Q (camera_module_cache_ram_94__4), 
         .QB (\$dummy [513]), .D (nx11803), .CLK (clk), .R (rst)) ;
    mux21_ni ix11804 (.Y (nx11803), .A0 (nx35432), .A1 (
             camera_module_cache_ram_94__4), .S0 (nx36674)) ;
    aoi22 ix26221 (.Y (nx26220), .A0 (camera_module_cache_ram_126__4), .A1 (
          nx36056), .B0 (camera_module_cache_ram_110__4), .B1 (nx36096)) ;
    dffr camera_module_cache_reg_ram_126__4 (.Q (camera_module_cache_ram_126__4)
         , .QB (\$dummy [514]), .D (nx11783), .CLK (clk), .R (rst)) ;
    mux21_ni ix11784 (.Y (nx11783), .A0 (nx35432), .A1 (
             camera_module_cache_ram_126__4), .S0 (nx36678)) ;
    dffr camera_module_cache_reg_ram_110__4 (.Q (camera_module_cache_ram_110__4)
         , .QB (\$dummy [515]), .D (nx11793), .CLK (clk), .R (rst)) ;
    mux21_ni ix11794 (.Y (nx11793), .A0 (nx35434), .A1 (
             camera_module_cache_ram_110__4), .S0 (nx36682)) ;
    nand04 ix14663 (.Y (nx14662), .A0 (nx26229), .A1 (nx26239), .A2 (nx26251), .A3 (
           nx26262)) ;
    aoi22 ix26230 (.Y (nx26229), .A0 (camera_module_cache_ram_142__4), .A1 (
          nx36136), .B0 (camera_module_cache_ram_158__4), .B1 (nx36176)) ;
    dffr camera_module_cache_reg_ram_142__4 (.Q (camera_module_cache_ram_142__4)
         , .QB (\$dummy [516]), .D (nx11773), .CLK (clk), .R (rst)) ;
    mux21_ni ix11774 (.Y (nx11773), .A0 (nx35434), .A1 (
             camera_module_cache_ram_142__4), .S0 (nx36686)) ;
    dffr camera_module_cache_reg_ram_158__4 (.Q (camera_module_cache_ram_158__4)
         , .QB (\$dummy [517]), .D (nx11763), .CLK (clk), .R (rst)) ;
    mux21_ni ix11764 (.Y (nx11763), .A0 (nx35434), .A1 (
             camera_module_cache_ram_158__4), .S0 (nx36690)) ;
    aoi22 ix26240 (.Y (nx26239), .A0 (camera_module_cache_ram_190__4), .A1 (
          nx36216), .B0 (camera_module_cache_ram_174__4), .B1 (nx36256)) ;
    dffr camera_module_cache_reg_ram_190__4 (.Q (camera_module_cache_ram_190__4)
         , .QB (\$dummy [518]), .D (nx11743), .CLK (clk), .R (rst)) ;
    mux21_ni ix11744 (.Y (nx11743), .A0 (nx35434), .A1 (
             camera_module_cache_ram_190__4), .S0 (nx36694)) ;
    dffr camera_module_cache_reg_ram_174__4 (.Q (camera_module_cache_ram_174__4)
         , .QB (\$dummy [519]), .D (nx11753), .CLK (clk), .R (rst)) ;
    mux21_ni ix11754 (.Y (nx11753), .A0 (nx35434), .A1 (
             camera_module_cache_ram_174__4), .S0 (nx36698)) ;
    aoi22 ix26252 (.Y (nx26251), .A0 (camera_module_cache_ram_206__4), .A1 (
          nx36296), .B0 (camera_module_cache_ram_222__4), .B1 (nx36336)) ;
    dffr camera_module_cache_reg_ram_206__4 (.Q (camera_module_cache_ram_206__4)
         , .QB (\$dummy [520]), .D (nx11733), .CLK (clk), .R (rst)) ;
    mux21_ni ix11734 (.Y (nx11733), .A0 (nx35434), .A1 (
             camera_module_cache_ram_206__4), .S0 (nx36702)) ;
    dffr camera_module_cache_reg_ram_222__4 (.Q (camera_module_cache_ram_222__4)
         , .QB (\$dummy [521]), .D (nx11723), .CLK (clk), .R (rst)) ;
    mux21_ni ix11724 (.Y (nx11723), .A0 (nx35434), .A1 (
             camera_module_cache_ram_222__4), .S0 (nx36706)) ;
    aoi22 ix26263 (.Y (nx26262), .A0 (camera_module_cache_ram_238__4), .A1 (
          nx36376), .B0 (camera_module_cache_ram_254__4), .B1 (nx36416)) ;
    dffr camera_module_cache_reg_ram_238__4 (.Q (camera_module_cache_ram_238__4)
         , .QB (\$dummy [522]), .D (nx11713), .CLK (clk), .R (rst)) ;
    mux21_ni ix11714 (.Y (nx11713), .A0 (nx35436), .A1 (
             camera_module_cache_ram_238__4), .S0 (nx36710)) ;
    dffr camera_module_cache_reg_ram_254__4 (.Q (camera_module_cache_ram_254__4)
         , .QB (\$dummy [523]), .D (nx11703), .CLK (clk), .R (rst)) ;
    mux21_ni ix11704 (.Y (nx11703), .A0 (nx35436), .A1 (
             camera_module_cache_ram_254__4), .S0 (nx36714)) ;
    oai21 ix26273 (.Y (nx26272), .A0 (nx14578), .A1 (nx14500), .B0 (nx36728)) ;
    nand04 ix14579 (.Y (nx14578), .A0 (nx26275), .A1 (nx26286), .A2 (nx26296), .A3 (
           nx26305)) ;
    aoi22 ix26276 (.Y (nx26275), .A0 (camera_module_cache_ram_15__4), .A1 (
          nx35818), .B0 (camera_module_cache_ram_31__4), .B1 (nx35858)) ;
    dffr camera_module_cache_reg_ram_15__4 (.Q (camera_module_cache_ram_15__4), 
         .QB (\$dummy [524]), .D (nx11693), .CLK (clk), .R (rst)) ;
    mux21_ni ix11694 (.Y (nx11693), .A0 (nx35436), .A1 (
             camera_module_cache_ram_15__4), .S0 (nx36718)) ;
    dffr camera_module_cache_reg_ram_31__4 (.Q (camera_module_cache_ram_31__4), 
         .QB (\$dummy [525]), .D (nx11683), .CLK (clk), .R (rst)) ;
    mux21_ni ix11684 (.Y (nx11683), .A0 (nx35436), .A1 (
             camera_module_cache_ram_31__4), .S0 (nx36732)) ;
    aoi22 ix26287 (.Y (nx26286), .A0 (camera_module_cache_ram_47__4), .A1 (
          nx35898), .B0 (camera_module_cache_ram_63__4), .B1 (nx35938)) ;
    dffr camera_module_cache_reg_ram_47__4 (.Q (camera_module_cache_ram_47__4), 
         .QB (\$dummy [526]), .D (nx11673), .CLK (clk), .R (rst)) ;
    mux21_ni ix11674 (.Y (nx11673), .A0 (nx35436), .A1 (
             camera_module_cache_ram_47__4), .S0 (nx36736)) ;
    dffr camera_module_cache_reg_ram_63__4 (.Q (camera_module_cache_ram_63__4), 
         .QB (\$dummy [527]), .D (nx11663), .CLK (clk), .R (rst)) ;
    mux21_ni ix11664 (.Y (nx11663), .A0 (nx35436), .A1 (
             camera_module_cache_ram_63__4), .S0 (nx36740)) ;
    aoi22 ix26297 (.Y (nx26296), .A0 (camera_module_cache_ram_79__4), .A1 (
          nx35978), .B0 (camera_module_cache_ram_95__4), .B1 (nx36018)) ;
    dffr camera_module_cache_reg_ram_79__4 (.Q (camera_module_cache_ram_79__4), 
         .QB (\$dummy [528]), .D (nx11653), .CLK (clk), .R (rst)) ;
    mux21_ni ix11654 (.Y (nx11653), .A0 (nx35436), .A1 (
             camera_module_cache_ram_79__4), .S0 (nx36744)) ;
    dffr camera_module_cache_reg_ram_95__4 (.Q (camera_module_cache_ram_95__4), 
         .QB (\$dummy [529]), .D (nx11643), .CLK (clk), .R (rst)) ;
    mux21_ni ix11644 (.Y (nx11643), .A0 (nx35438), .A1 (
             camera_module_cache_ram_95__4), .S0 (nx36748)) ;
    aoi22 ix26306 (.Y (nx26305), .A0 (camera_module_cache_ram_127__4), .A1 (
          nx36058), .B0 (camera_module_cache_ram_111__4), .B1 (nx36098)) ;
    dffr camera_module_cache_reg_ram_127__4 (.Q (camera_module_cache_ram_127__4)
         , .QB (\$dummy [530]), .D (nx11623), .CLK (clk), .R (rst)) ;
    mux21_ni ix11624 (.Y (nx11623), .A0 (nx35438), .A1 (
             camera_module_cache_ram_127__4), .S0 (nx36752)) ;
    dffr camera_module_cache_reg_ram_111__4 (.Q (camera_module_cache_ram_111__4)
         , .QB (\$dummy [531]), .D (nx11633), .CLK (clk), .R (rst)) ;
    mux21_ni ix11634 (.Y (nx11633), .A0 (nx35438), .A1 (
             camera_module_cache_ram_111__4), .S0 (nx36756)) ;
    nand04 ix14501 (.Y (nx14500), .A0 (nx26315), .A1 (nx26327), .A2 (nx26339), .A3 (
           nx26349)) ;
    aoi22 ix26316 (.Y (nx26315), .A0 (camera_module_cache_ram_143__4), .A1 (
          nx36138), .B0 (camera_module_cache_ram_159__4), .B1 (nx36178)) ;
    dffr camera_module_cache_reg_ram_143__4 (.Q (camera_module_cache_ram_143__4)
         , .QB (\$dummy [532]), .D (nx11613), .CLK (clk), .R (rst)) ;
    mux21_ni ix11614 (.Y (nx11613), .A0 (nx35438), .A1 (
             camera_module_cache_ram_143__4), .S0 (nx36760)) ;
    dffr camera_module_cache_reg_ram_159__4 (.Q (camera_module_cache_ram_159__4)
         , .QB (\$dummy [533]), .D (nx11603), .CLK (clk), .R (rst)) ;
    mux21_ni ix11604 (.Y (nx11603), .A0 (nx35438), .A1 (
             camera_module_cache_ram_159__4), .S0 (nx36764)) ;
    aoi22 ix26328 (.Y (nx26327), .A0 (camera_module_cache_ram_191__4), .A1 (
          nx36218), .B0 (camera_module_cache_ram_175__4), .B1 (nx36258)) ;
    dffr camera_module_cache_reg_ram_191__4 (.Q (camera_module_cache_ram_191__4)
         , .QB (\$dummy [534]), .D (nx11583), .CLK (clk), .R (rst)) ;
    mux21_ni ix11584 (.Y (nx11583), .A0 (nx35438), .A1 (
             camera_module_cache_ram_191__4), .S0 (nx36768)) ;
    dffr camera_module_cache_reg_ram_175__4 (.Q (camera_module_cache_ram_175__4)
         , .QB (\$dummy [535]), .D (nx11593), .CLK (clk), .R (rst)) ;
    mux21_ni ix11594 (.Y (nx11593), .A0 (nx35438), .A1 (
             camera_module_cache_ram_175__4), .S0 (nx36772)) ;
    aoi22 ix26340 (.Y (nx26339), .A0 (camera_module_cache_ram_207__4), .A1 (
          nx36298), .B0 (camera_module_cache_ram_223__4), .B1 (nx36338)) ;
    dffr camera_module_cache_reg_ram_207__4 (.Q (camera_module_cache_ram_207__4)
         , .QB (\$dummy [536]), .D (nx11573), .CLK (clk), .R (rst)) ;
    mux21_ni ix11574 (.Y (nx11573), .A0 (nx35440), .A1 (
             camera_module_cache_ram_207__4), .S0 (nx36776)) ;
    dffr camera_module_cache_reg_ram_223__4 (.Q (camera_module_cache_ram_223__4)
         , .QB (\$dummy [537]), .D (nx11563), .CLK (clk), .R (rst)) ;
    mux21_ni ix11564 (.Y (nx11563), .A0 (nx35440), .A1 (
             camera_module_cache_ram_223__4), .S0 (nx36780)) ;
    aoi22 ix26350 (.Y (nx26349), .A0 (camera_module_cache_ram_239__4), .A1 (
          nx36378), .B0 (camera_module_cache_ram_255__4), .B1 (nx36418)) ;
    dffr camera_module_cache_reg_ram_239__4 (.Q (camera_module_cache_ram_239__4)
         , .QB (\$dummy [538]), .D (nx11553), .CLK (clk), .R (rst)) ;
    mux21_ni ix11554 (.Y (nx11553), .A0 (nx35440), .A1 (
             camera_module_cache_ram_239__4), .S0 (nx36784)) ;
    dffr camera_module_cache_reg_ram_255__4 (.Q (camera_module_cache_ram_255__4)
         , .QB (\$dummy [539]), .D (nx11543), .CLK (clk), .R (rst)) ;
    mux21_ni ix11544 (.Y (nx11543), .A0 (nx35440), .A1 (
             camera_module_cache_ram_255__4), .S0 (nx36788)) ;
    oai22 ix14303 (.Y (nx14302), .A0 (nx26363), .A1 (nx29959), .B0 (nx31098), .B1 (
          nx14278)) ;
    aoi22 ix26364 (.Y (nx26363), .A0 (camera_module_algo_module_pixel_value_2), 
          .A1 (nx26370), .B0 (nx8754), .B1 (nx11520)) ;
    dff camera_module_algo_module_pixel_reg_reg_q_2 (.Q (
        camera_module_algo_module_pixel_value_2), .QB (\$dummy [540]), .D (
        nx8963), .CLK (clk)) ;
    mux21_ni ix8964 (.Y (nx8963), .A0 (nx11512), .A1 (
             camera_module_algo_module_pixel_value_2), .S0 (nx37152)) ;
    mux21_ni ix26371 (.Y (nx26370), .A0 (nx26372), .A1 (nx35674), .S0 (nx36792)
             ) ;
    nor04 ix26373 (.Y (nx26372), .A0 (nx11492), .A1 (nx10838), .A2 (nx10182), .A3 (
          nx9528)) ;
    nand04 ix11493 (.Y (nx11492), .A0 (nx26375), .A1 (nx26521), .A2 (nx26600), .A3 (
           nx26680)) ;
    oai21 ix26376 (.Y (nx26375), .A0 (nx11482), .A1 (nx11404), .B0 (nx36448)) ;
    nand04 ix11483 (.Y (nx11482), .A0 (nx26379), .A1 (nx26444), .A2 (nx26453), .A3 (
           nx26463)) ;
    aoi22 ix26380 (.Y (nx26379), .A0 (camera_module_cache_ram_0__2), .A1 (
          nx35818), .B0 (camera_module_cache_ram_16__2), .B1 (nx35858)) ;
    dffr camera_module_cache_reg_ram_0__2 (.Q (camera_module_cache_ram_0__2), .QB (
         \$dummy [541]), .D (nx8953), .CLK (clk), .R (rst)) ;
    mux21_ni ix8954 (.Y (nx8953), .A0 (camera_module_cache_ram_0__2), .A1 (
             nx35216), .S0 (nx35134)) ;
    oai221 ix8875 (.Y (nx8874), .A0 (nx34074), .A1 (nx26385), .B0 (nx26411), .B1 (
           nx35712), .C0 (nx26415)) ;
    tri01 nvm_module_tri_dataout_122 (.Y (nvm_data_122), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_114 (.Y (nvm_data_114), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_106 (.Y (nvm_data_106), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_98 (.Y (nvm_data_98), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_90 (.Y (nvm_data_90), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_82 (.Y (nvm_data_82), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_74 (.Y (nvm_data_74), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_66 (.Y (nvm_data_66), .A (nx22549), .E (
          nvm_module_GND0)) ;
    inv01 ix26412 (.Y (nx26411), .A (nvm_data_2)) ;
    tri01 nvm_module_tri_dataout_2 (.Y (nvm_data_2), .A (nx22549), .E (
          nvm_module_GND0)) ;
    nand02 ix26416 (.Y (nx26415), .A0 (nx34074), .A1 (nx8808)) ;
    tri01 nvm_module_tri_dataout_58 (.Y (nvm_data_58), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_50 (.Y (nvm_data_50), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_42 (.Y (nvm_data_42), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_34 (.Y (nvm_data_34), .A (nx22549), .E (
          nvm_module_GND0)) ;
    oai22 ix8777 (.Y (nx8776), .A0 (nx34102), .A1 (nx26429), .B0 (nx34084), .B1 (
          nx26435)) ;
    tri01 nvm_module_tri_dataout_26 (.Y (nvm_data_26), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_18 (.Y (nvm_data_18), .A (nx22549), .E (
          nvm_module_GND0)) ;
    nand02 ix26436 (.Y (nx26435), .A0 (nvm_data_10), .A1 (nx34102)) ;
    tri01 nvm_module_tri_dataout_10 (.Y (nvm_data_10), .A (nx22549), .E (
          nvm_module_GND0)) ;
    dffr camera_module_cache_reg_ram_16__2 (.Q (camera_module_cache_ram_16__2), 
         .QB (\$dummy [542]), .D (nx8943), .CLK (clk), .R (rst)) ;
    mux21_ni ix8944 (.Y (nx8943), .A0 (camera_module_cache_ram_16__2), .A1 (
             nx35216), .S0 (nx35130)) ;
    aoi22 ix26445 (.Y (nx26444), .A0 (camera_module_cache_ram_32__2), .A1 (
          nx35898), .B0 (camera_module_cache_ram_48__2), .B1 (nx35938)) ;
    dffr camera_module_cache_reg_ram_32__2 (.Q (camera_module_cache_ram_32__2), 
         .QB (\$dummy [543]), .D (nx8933), .CLK (clk), .R (rst)) ;
    mux21_ni ix8934 (.Y (nx8933), .A0 (camera_module_cache_ram_32__2), .A1 (
             nx35216), .S0 (nx35126)) ;
    dffr camera_module_cache_reg_ram_48__2 (.Q (camera_module_cache_ram_48__2), 
         .QB (\$dummy [544]), .D (nx8923), .CLK (clk), .R (rst)) ;
    mux21_ni ix8924 (.Y (nx8923), .A0 (camera_module_cache_ram_48__2), .A1 (
             nx35216), .S0 (nx35122)) ;
    aoi22 ix26454 (.Y (nx26453), .A0 (camera_module_cache_ram_64__2), .A1 (
          nx35978), .B0 (camera_module_cache_ram_80__2), .B1 (nx36018)) ;
    dffr camera_module_cache_reg_ram_64__2 (.Q (camera_module_cache_ram_64__2), 
         .QB (\$dummy [545]), .D (nx8913), .CLK (clk), .R (rst)) ;
    mux21_ni ix8914 (.Y (nx8913), .A0 (camera_module_cache_ram_64__2), .A1 (
             nx35216), .S0 (nx35118)) ;
    dffr camera_module_cache_reg_ram_80__2 (.Q (camera_module_cache_ram_80__2), 
         .QB (\$dummy [546]), .D (nx8903), .CLK (clk), .R (rst)) ;
    mux21_ni ix8904 (.Y (nx8903), .A0 (camera_module_cache_ram_80__2), .A1 (
             nx35216), .S0 (nx35114)) ;
    aoi22 ix26464 (.Y (nx26463), .A0 (camera_module_cache_ram_112__2), .A1 (
          nx36058), .B0 (camera_module_cache_ram_96__2), .B1 (nx36098)) ;
    dffr camera_module_cache_reg_ram_112__2 (.Q (camera_module_cache_ram_112__2)
         , .QB (\$dummy [547]), .D (nx8883), .CLK (clk), .R (rst)) ;
    mux21_ni ix8884 (.Y (nx8883), .A0 (camera_module_cache_ram_112__2), .A1 (
             nx35216), .S0 (nx35106)) ;
    dffr camera_module_cache_reg_ram_96__2 (.Q (camera_module_cache_ram_96__2), 
         .QB (\$dummy [548]), .D (nx8893), .CLK (clk), .R (rst)) ;
    mux21_ni ix8894 (.Y (nx8893), .A0 (camera_module_cache_ram_96__2), .A1 (
             nx35218), .S0 (nx35110)) ;
    nand04 ix11405 (.Y (nx11404), .A0 (nx26475), .A1 (nx26487), .A2 (nx26497), .A3 (
           nx26508)) ;
    aoi22 ix26476 (.Y (nx26475), .A0 (camera_module_cache_ram_128__2), .A1 (
          nx36138), .B0 (camera_module_cache_ram_144__2), .B1 (nx36178)) ;
    dffr camera_module_cache_reg_ram_128__2 (.Q (camera_module_cache_ram_128__2)
         , .QB (\$dummy [549]), .D (nx8873), .CLK (clk), .R (rst)) ;
    mux21_ni ix8874 (.Y (nx8873), .A0 (camera_module_cache_ram_128__2), .A1 (
             nx35218), .S0 (nx35102)) ;
    dffr camera_module_cache_reg_ram_144__2 (.Q (camera_module_cache_ram_144__2)
         , .QB (\$dummy [550]), .D (nx8863), .CLK (clk), .R (rst)) ;
    mux21_ni ix8864 (.Y (nx8863), .A0 (camera_module_cache_ram_144__2), .A1 (
             nx35218), .S0 (nx35098)) ;
    aoi22 ix26488 (.Y (nx26487), .A0 (camera_module_cache_ram_176__2), .A1 (
          nx36218), .B0 (camera_module_cache_ram_160__2), .B1 (nx36258)) ;
    dffr camera_module_cache_reg_ram_176__2 (.Q (camera_module_cache_ram_176__2)
         , .QB (\$dummy [551]), .D (nx8843), .CLK (clk), .R (rst)) ;
    mux21_ni ix8844 (.Y (nx8843), .A0 (camera_module_cache_ram_176__2), .A1 (
             nx35218), .S0 (nx35090)) ;
    dffr camera_module_cache_reg_ram_160__2 (.Q (camera_module_cache_ram_160__2)
         , .QB (\$dummy [552]), .D (nx8853), .CLK (clk), .R (rst)) ;
    mux21_ni ix8854 (.Y (nx8853), .A0 (camera_module_cache_ram_160__2), .A1 (
             nx35218), .S0 (nx35094)) ;
    aoi22 ix26498 (.Y (nx26497), .A0 (camera_module_cache_ram_192__2), .A1 (
          nx36298), .B0 (camera_module_cache_ram_208__2), .B1 (nx36338)) ;
    dffr camera_module_cache_reg_ram_192__2 (.Q (camera_module_cache_ram_192__2)
         , .QB (\$dummy [553]), .D (nx8833), .CLK (clk), .R (rst)) ;
    mux21_ni ix8834 (.Y (nx8833), .A0 (camera_module_cache_ram_192__2), .A1 (
             nx35218), .S0 (nx35086)) ;
    dffr camera_module_cache_reg_ram_208__2 (.Q (camera_module_cache_ram_208__2)
         , .QB (\$dummy [554]), .D (nx8823), .CLK (clk), .R (rst)) ;
    mux21_ni ix8824 (.Y (nx8823), .A0 (camera_module_cache_ram_208__2), .A1 (
             nx35218), .S0 (nx35082)) ;
    aoi22 ix26510 (.Y (nx26508), .A0 (camera_module_cache_ram_224__2), .A1 (
          nx36378), .B0 (camera_module_cache_ram_240__2), .B1 (nx36418)) ;
    dffr camera_module_cache_reg_ram_224__2 (.Q (camera_module_cache_ram_224__2)
         , .QB (\$dummy [555]), .D (nx8813), .CLK (clk), .R (rst)) ;
    mux21_ni ix8814 (.Y (nx8813), .A0 (camera_module_cache_ram_224__2), .A1 (
             nx35220), .S0 (nx35078)) ;
    dffr camera_module_cache_reg_ram_240__2 (.Q (camera_module_cache_ram_240__2)
         , .QB (\$dummy [556]), .D (nx8803), .CLK (clk), .R (rst)) ;
    mux21_ni ix8804 (.Y (nx8803), .A0 (camera_module_cache_ram_240__2), .A1 (
             nx35220), .S0 (nx35074)) ;
    oai21 ix26522 (.Y (nx26521), .A0 (nx11320), .A1 (nx11242), .B0 (nx36452)) ;
    nand04 ix11321 (.Y (nx11320), .A0 (nx26525), .A1 (nx26536), .A2 (nx26545), .A3 (
           nx26554)) ;
    aoi22 ix26526 (.Y (nx26525), .A0 (camera_module_cache_ram_1__2), .A1 (
          nx35818), .B0 (camera_module_cache_ram_17__2), .B1 (nx35858)) ;
    dffr camera_module_cache_reg_ram_1__2 (.Q (camera_module_cache_ram_1__2), .QB (
         \$dummy [557]), .D (nx8793), .CLK (clk), .R (rst)) ;
    mux21_ni ix8794 (.Y (nx8793), .A0 (camera_module_cache_ram_1__2), .A1 (
             nx35220), .S0 (nx35064)) ;
    dffr camera_module_cache_reg_ram_17__2 (.Q (camera_module_cache_ram_17__2), 
         .QB (\$dummy [558]), .D (nx8783), .CLK (clk), .R (rst)) ;
    mux21_ni ix8784 (.Y (nx8783), .A0 (camera_module_cache_ram_17__2), .A1 (
             nx35220), .S0 (nx35060)) ;
    aoi22 ix26537 (.Y (nx26536), .A0 (camera_module_cache_ram_33__2), .A1 (
          nx35898), .B0 (camera_module_cache_ram_49__2), .B1 (nx35938)) ;
    dffr camera_module_cache_reg_ram_33__2 (.Q (camera_module_cache_ram_33__2), 
         .QB (\$dummy [559]), .D (nx8773), .CLK (clk), .R (rst)) ;
    mux21_ni ix8774 (.Y (nx8773), .A0 (camera_module_cache_ram_33__2), .A1 (
             nx35220), .S0 (nx35056)) ;
    dffr camera_module_cache_reg_ram_49__2 (.Q (camera_module_cache_ram_49__2), 
         .QB (\$dummy [560]), .D (nx8763), .CLK (clk), .R (rst)) ;
    mux21_ni ix8764 (.Y (nx8763), .A0 (camera_module_cache_ram_49__2), .A1 (
             nx35220), .S0 (nx35052)) ;
    aoi22 ix26546 (.Y (nx26545), .A0 (camera_module_cache_ram_65__2), .A1 (
          nx35978), .B0 (camera_module_cache_ram_81__2), .B1 (nx36018)) ;
    dffr camera_module_cache_reg_ram_65__2 (.Q (camera_module_cache_ram_65__2), 
         .QB (\$dummy [561]), .D (nx8753), .CLK (clk), .R (rst)) ;
    mux21_ni ix8754 (.Y (nx8753), .A0 (camera_module_cache_ram_65__2), .A1 (
             nx35220), .S0 (nx35048)) ;
    dffr camera_module_cache_reg_ram_81__2 (.Q (camera_module_cache_ram_81__2), 
         .QB (\$dummy [562]), .D (nx8743), .CLK (clk), .R (rst)) ;
    mux21_ni ix8744 (.Y (nx8743), .A0 (camera_module_cache_ram_81__2), .A1 (
             nx35222), .S0 (nx35044)) ;
    aoi22 ix26555 (.Y (nx26554), .A0 (camera_module_cache_ram_113__2), .A1 (
          nx36058), .B0 (camera_module_cache_ram_97__2), .B1 (nx36098)) ;
    dffr camera_module_cache_reg_ram_113__2 (.Q (camera_module_cache_ram_113__2)
         , .QB (\$dummy [563]), .D (nx8723), .CLK (clk), .R (rst)) ;
    mux21_ni ix8724 (.Y (nx8723), .A0 (camera_module_cache_ram_113__2), .A1 (
             nx35222), .S0 (nx35036)) ;
    dffr camera_module_cache_reg_ram_97__2 (.Q (camera_module_cache_ram_97__2), 
         .QB (\$dummy [564]), .D (nx8733), .CLK (clk), .R (rst)) ;
    mux21_ni ix8734 (.Y (nx8733), .A0 (camera_module_cache_ram_97__2), .A1 (
             nx35222), .S0 (nx35040)) ;
    nand04 ix11243 (.Y (nx11242), .A0 (nx26563), .A1 (nx26573), .A2 (nx26582), .A3 (
           nx26590)) ;
    aoi22 ix26564 (.Y (nx26563), .A0 (camera_module_cache_ram_129__2), .A1 (
          nx36138), .B0 (camera_module_cache_ram_145__2), .B1 (nx36178)) ;
    dffr camera_module_cache_reg_ram_129__2 (.Q (camera_module_cache_ram_129__2)
         , .QB (\$dummy [565]), .D (nx8713), .CLK (clk), .R (rst)) ;
    mux21_ni ix8714 (.Y (nx8713), .A0 (camera_module_cache_ram_129__2), .A1 (
             nx35222), .S0 (nx35032)) ;
    dffr camera_module_cache_reg_ram_145__2 (.Q (camera_module_cache_ram_145__2)
         , .QB (\$dummy [566]), .D (nx8703), .CLK (clk), .R (rst)) ;
    mux21_ni ix8704 (.Y (nx8703), .A0 (camera_module_cache_ram_145__2), .A1 (
             nx35222), .S0 (nx35028)) ;
    aoi22 ix26574 (.Y (nx26573), .A0 (camera_module_cache_ram_177__2), .A1 (
          nx36218), .B0 (camera_module_cache_ram_161__2), .B1 (nx36258)) ;
    dffr camera_module_cache_reg_ram_177__2 (.Q (camera_module_cache_ram_177__2)
         , .QB (\$dummy [567]), .D (nx8683), .CLK (clk), .R (rst)) ;
    mux21_ni ix8684 (.Y (nx8683), .A0 (camera_module_cache_ram_177__2), .A1 (
             nx35222), .S0 (nx35020)) ;
    dffr camera_module_cache_reg_ram_161__2 (.Q (camera_module_cache_ram_161__2)
         , .QB (\$dummy [568]), .D (nx8693), .CLK (clk), .R (rst)) ;
    mux21_ni ix8694 (.Y (nx8693), .A0 (camera_module_cache_ram_161__2), .A1 (
             nx35222), .S0 (nx35024)) ;
    aoi22 ix26583 (.Y (nx26582), .A0 (camera_module_cache_ram_193__2), .A1 (
          nx36298), .B0 (camera_module_cache_ram_209__2), .B1 (nx36338)) ;
    dffr camera_module_cache_reg_ram_193__2 (.Q (camera_module_cache_ram_193__2)
         , .QB (\$dummy [569]), .D (nx8673), .CLK (clk), .R (rst)) ;
    mux21_ni ix8674 (.Y (nx8673), .A0 (camera_module_cache_ram_193__2), .A1 (
             nx35224), .S0 (nx35016)) ;
    dffr camera_module_cache_reg_ram_209__2 (.Q (camera_module_cache_ram_209__2)
         , .QB (\$dummy [570]), .D (nx8663), .CLK (clk), .R (rst)) ;
    mux21_ni ix8664 (.Y (nx8663), .A0 (camera_module_cache_ram_209__2), .A1 (
             nx35224), .S0 (nx35012)) ;
    aoi22 ix26591 (.Y (nx26590), .A0 (camera_module_cache_ram_225__2), .A1 (
          nx36378), .B0 (camera_module_cache_ram_241__2), .B1 (nx36418)) ;
    dffr camera_module_cache_reg_ram_225__2 (.Q (camera_module_cache_ram_225__2)
         , .QB (\$dummy [571]), .D (nx8653), .CLK (clk), .R (rst)) ;
    mux21_ni ix8654 (.Y (nx8653), .A0 (camera_module_cache_ram_225__2), .A1 (
             nx35224), .S0 (nx35008)) ;
    dffr camera_module_cache_reg_ram_241__2 (.Q (camera_module_cache_ram_241__2)
         , .QB (\$dummy [572]), .D (nx8643), .CLK (clk), .R (rst)) ;
    mux21_ni ix8644 (.Y (nx8643), .A0 (camera_module_cache_ram_241__2), .A1 (
             nx35224), .S0 (nx35004)) ;
    oai21 ix26601 (.Y (nx26600), .A0 (nx11156), .A1 (nx11078), .B0 (nx36456)) ;
    nand04 ix11157 (.Y (nx11156), .A0 (nx26603), .A1 (nx26614), .A2 (nx26622), .A3 (
           nx26632)) ;
    aoi22 ix26604 (.Y (nx26603), .A0 (camera_module_cache_ram_2__2), .A1 (
          nx35818), .B0 (camera_module_cache_ram_18__2), .B1 (nx35858)) ;
    dffr camera_module_cache_reg_ram_2__2 (.Q (camera_module_cache_ram_2__2), .QB (
         \$dummy [573]), .D (nx8633), .CLK (clk), .R (rst)) ;
    mux21_ni ix8634 (.Y (nx8633), .A0 (camera_module_cache_ram_2__2), .A1 (
             nx35224), .S0 (nx34994)) ;
    dffr camera_module_cache_reg_ram_18__2 (.Q (camera_module_cache_ram_18__2), 
         .QB (\$dummy [574]), .D (nx8623), .CLK (clk), .R (rst)) ;
    mux21_ni ix8624 (.Y (nx8623), .A0 (camera_module_cache_ram_18__2), .A1 (
             nx35224), .S0 (nx34990)) ;
    aoi22 ix26615 (.Y (nx26614), .A0 (camera_module_cache_ram_34__2), .A1 (
          nx35898), .B0 (camera_module_cache_ram_50__2), .B1 (nx35938)) ;
    dffr camera_module_cache_reg_ram_34__2 (.Q (camera_module_cache_ram_34__2), 
         .QB (\$dummy [575]), .D (nx8613), .CLK (clk), .R (rst)) ;
    mux21_ni ix8614 (.Y (nx8613), .A0 (camera_module_cache_ram_34__2), .A1 (
             nx35224), .S0 (nx34986)) ;
    dffr camera_module_cache_reg_ram_50__2 (.Q (camera_module_cache_ram_50__2), 
         .QB (\$dummy [576]), .D (nx8603), .CLK (clk), .R (rst)) ;
    mux21_ni ix8604 (.Y (nx8603), .A0 (camera_module_cache_ram_50__2), .A1 (
             nx35226), .S0 (nx34982)) ;
    aoi22 ix26623 (.Y (nx26622), .A0 (camera_module_cache_ram_66__2), .A1 (
          nx35978), .B0 (camera_module_cache_ram_82__2), .B1 (nx36018)) ;
    dffr camera_module_cache_reg_ram_66__2 (.Q (camera_module_cache_ram_66__2), 
         .QB (\$dummy [577]), .D (nx8593), .CLK (clk), .R (rst)) ;
    mux21_ni ix8594 (.Y (nx8593), .A0 (camera_module_cache_ram_66__2), .A1 (
             nx35226), .S0 (nx34978)) ;
    dffr camera_module_cache_reg_ram_82__2 (.Q (camera_module_cache_ram_82__2), 
         .QB (\$dummy [578]), .D (nx8583), .CLK (clk), .R (rst)) ;
    mux21_ni ix8584 (.Y (nx8583), .A0 (camera_module_cache_ram_82__2), .A1 (
             nx35226), .S0 (nx34974)) ;
    aoi22 ix26633 (.Y (nx26632), .A0 (camera_module_cache_ram_114__2), .A1 (
          nx36058), .B0 (camera_module_cache_ram_98__2), .B1 (nx36098)) ;
    dffr camera_module_cache_reg_ram_114__2 (.Q (camera_module_cache_ram_114__2)
         , .QB (\$dummy [579]), .D (nx8563), .CLK (clk), .R (rst)) ;
    mux21_ni ix8564 (.Y (nx8563), .A0 (camera_module_cache_ram_114__2), .A1 (
             nx35226), .S0 (nx34966)) ;
    dffr camera_module_cache_reg_ram_98__2 (.Q (camera_module_cache_ram_98__2), 
         .QB (\$dummy [580]), .D (nx8573), .CLK (clk), .R (rst)) ;
    mux21_ni ix8574 (.Y (nx8573), .A0 (camera_module_cache_ram_98__2), .A1 (
             nx35226), .S0 (nx34970)) ;
    nand04 ix11079 (.Y (nx11078), .A0 (nx26643), .A1 (nx26653), .A2 (nx26662), .A3 (
           nx26670)) ;
    aoi22 ix26644 (.Y (nx26643), .A0 (camera_module_cache_ram_130__2), .A1 (
          nx36138), .B0 (camera_module_cache_ram_146__2), .B1 (nx36178)) ;
    dffr camera_module_cache_reg_ram_130__2 (.Q (camera_module_cache_ram_130__2)
         , .QB (\$dummy [581]), .D (nx8553), .CLK (clk), .R (rst)) ;
    mux21_ni ix8554 (.Y (nx8553), .A0 (camera_module_cache_ram_130__2), .A1 (
             nx35226), .S0 (nx34962)) ;
    dffr camera_module_cache_reg_ram_146__2 (.Q (camera_module_cache_ram_146__2)
         , .QB (\$dummy [582]), .D (nx8543), .CLK (clk), .R (rst)) ;
    mux21_ni ix8544 (.Y (nx8543), .A0 (camera_module_cache_ram_146__2), .A1 (
             nx35226), .S0 (nx34958)) ;
    aoi22 ix26654 (.Y (nx26653), .A0 (camera_module_cache_ram_178__2), .A1 (
          nx36218), .B0 (camera_module_cache_ram_162__2), .B1 (nx36258)) ;
    dffr camera_module_cache_reg_ram_178__2 (.Q (camera_module_cache_ram_178__2)
         , .QB (\$dummy [583]), .D (nx8523), .CLK (clk), .R (rst)) ;
    mux21_ni ix8524 (.Y (nx8523), .A0 (camera_module_cache_ram_178__2), .A1 (
             nx35228), .S0 (nx34950)) ;
    dffr camera_module_cache_reg_ram_162__2 (.Q (camera_module_cache_ram_162__2)
         , .QB (\$dummy [584]), .D (nx8533), .CLK (clk), .R (rst)) ;
    mux21_ni ix8534 (.Y (nx8533), .A0 (camera_module_cache_ram_162__2), .A1 (
             nx35228), .S0 (nx34954)) ;
    aoi22 ix26663 (.Y (nx26662), .A0 (camera_module_cache_ram_194__2), .A1 (
          nx36298), .B0 (camera_module_cache_ram_210__2), .B1 (nx36338)) ;
    dffr camera_module_cache_reg_ram_194__2 (.Q (camera_module_cache_ram_194__2)
         , .QB (\$dummy [585]), .D (nx8513), .CLK (clk), .R (rst)) ;
    mux21_ni ix8514 (.Y (nx8513), .A0 (camera_module_cache_ram_194__2), .A1 (
             nx35228), .S0 (nx34946)) ;
    dffr camera_module_cache_reg_ram_210__2 (.Q (camera_module_cache_ram_210__2)
         , .QB (\$dummy [586]), .D (nx8503), .CLK (clk), .R (rst)) ;
    mux21_ni ix8504 (.Y (nx8503), .A0 (camera_module_cache_ram_210__2), .A1 (
             nx35228), .S0 (nx34942)) ;
    aoi22 ix26671 (.Y (nx26670), .A0 (camera_module_cache_ram_226__2), .A1 (
          nx36378), .B0 (camera_module_cache_ram_242__2), .B1 (nx36418)) ;
    dffr camera_module_cache_reg_ram_226__2 (.Q (camera_module_cache_ram_226__2)
         , .QB (\$dummy [587]), .D (nx8493), .CLK (clk), .R (rst)) ;
    mux21_ni ix8494 (.Y (nx8493), .A0 (camera_module_cache_ram_226__2), .A1 (
             nx35228), .S0 (nx34938)) ;
    dffr camera_module_cache_reg_ram_242__2 (.Q (camera_module_cache_ram_242__2)
         , .QB (\$dummy [588]), .D (nx8483), .CLK (clk), .R (rst)) ;
    mux21_ni ix8484 (.Y (nx8483), .A0 (camera_module_cache_ram_242__2), .A1 (
             nx35228), .S0 (nx34934)) ;
    oai21 ix26681 (.Y (nx26680), .A0 (nx10994), .A1 (nx10916), .B0 (nx36460)) ;
    nand04 ix10995 (.Y (nx10994), .A0 (nx26683), .A1 (nx26694), .A2 (nx26702), .A3 (
           nx26712)) ;
    aoi22 ix26684 (.Y (nx26683), .A0 (camera_module_cache_ram_3__2), .A1 (
          nx35818), .B0 (camera_module_cache_ram_19__2), .B1 (nx35858)) ;
    dffr camera_module_cache_reg_ram_3__2 (.Q (camera_module_cache_ram_3__2), .QB (
         \$dummy [589]), .D (nx8473), .CLK (clk), .R (rst)) ;
    mux21_ni ix8474 (.Y (nx8473), .A0 (camera_module_cache_ram_3__2), .A1 (
             nx35228), .S0 (nx34924)) ;
    dffr camera_module_cache_reg_ram_19__2 (.Q (camera_module_cache_ram_19__2), 
         .QB (\$dummy [590]), .D (nx8463), .CLK (clk), .R (rst)) ;
    mux21_ni ix8464 (.Y (nx8463), .A0 (camera_module_cache_ram_19__2), .A1 (
             nx35230), .S0 (nx34920)) ;
    aoi22 ix26695 (.Y (nx26694), .A0 (camera_module_cache_ram_35__2), .A1 (
          nx35898), .B0 (camera_module_cache_ram_51__2), .B1 (nx35938)) ;
    dffr camera_module_cache_reg_ram_35__2 (.Q (camera_module_cache_ram_35__2), 
         .QB (\$dummy [591]), .D (nx8453), .CLK (clk), .R (rst)) ;
    mux21_ni ix8454 (.Y (nx8453), .A0 (camera_module_cache_ram_35__2), .A1 (
             nx35230), .S0 (nx34916)) ;
    dffr camera_module_cache_reg_ram_51__2 (.Q (camera_module_cache_ram_51__2), 
         .QB (\$dummy [592]), .D (nx8443), .CLK (clk), .R (rst)) ;
    mux21_ni ix8444 (.Y (nx8443), .A0 (camera_module_cache_ram_51__2), .A1 (
             nx35230), .S0 (nx34912)) ;
    aoi22 ix26703 (.Y (nx26702), .A0 (camera_module_cache_ram_67__2), .A1 (
          nx35978), .B0 (camera_module_cache_ram_83__2), .B1 (nx36018)) ;
    dffr camera_module_cache_reg_ram_67__2 (.Q (camera_module_cache_ram_67__2), 
         .QB (\$dummy [593]), .D (nx8433), .CLK (clk), .R (rst)) ;
    mux21_ni ix8434 (.Y (nx8433), .A0 (camera_module_cache_ram_67__2), .A1 (
             nx35230), .S0 (nx34908)) ;
    dffr camera_module_cache_reg_ram_83__2 (.Q (camera_module_cache_ram_83__2), 
         .QB (\$dummy [594]), .D (nx8423), .CLK (clk), .R (rst)) ;
    mux21_ni ix8424 (.Y (nx8423), .A0 (camera_module_cache_ram_83__2), .A1 (
             nx35230), .S0 (nx34904)) ;
    aoi22 ix26713 (.Y (nx26712), .A0 (camera_module_cache_ram_115__2), .A1 (
          nx36058), .B0 (camera_module_cache_ram_99__2), .B1 (nx36098)) ;
    dffr camera_module_cache_reg_ram_115__2 (.Q (camera_module_cache_ram_115__2)
         , .QB (\$dummy [595]), .D (nx8403), .CLK (clk), .R (rst)) ;
    mux21_ni ix8404 (.Y (nx8403), .A0 (camera_module_cache_ram_115__2), .A1 (
             nx35230), .S0 (nx34896)) ;
    dffr camera_module_cache_reg_ram_99__2 (.Q (camera_module_cache_ram_99__2), 
         .QB (\$dummy [596]), .D (nx8413), .CLK (clk), .R (rst)) ;
    mux21_ni ix8414 (.Y (nx8413), .A0 (camera_module_cache_ram_99__2), .A1 (
             nx35230), .S0 (nx34900)) ;
    nand04 ix10917 (.Y (nx10916), .A0 (nx26723), .A1 (nx26733), .A2 (nx26742), .A3 (
           nx26750)) ;
    aoi22 ix26724 (.Y (nx26723), .A0 (camera_module_cache_ram_131__2), .A1 (
          nx36138), .B0 (camera_module_cache_ram_147__2), .B1 (nx36178)) ;
    dffr camera_module_cache_reg_ram_131__2 (.Q (camera_module_cache_ram_131__2)
         , .QB (\$dummy [597]), .D (nx8393), .CLK (clk), .R (rst)) ;
    mux21_ni ix8394 (.Y (nx8393), .A0 (camera_module_cache_ram_131__2), .A1 (
             nx35232), .S0 (nx34892)) ;
    dffr camera_module_cache_reg_ram_147__2 (.Q (camera_module_cache_ram_147__2)
         , .QB (\$dummy [598]), .D (nx8383), .CLK (clk), .R (rst)) ;
    mux21_ni ix8384 (.Y (nx8383), .A0 (camera_module_cache_ram_147__2), .A1 (
             nx35232), .S0 (nx34888)) ;
    aoi22 ix26734 (.Y (nx26733), .A0 (camera_module_cache_ram_179__2), .A1 (
          nx36218), .B0 (camera_module_cache_ram_163__2), .B1 (nx36258)) ;
    dffr camera_module_cache_reg_ram_179__2 (.Q (camera_module_cache_ram_179__2)
         , .QB (\$dummy [599]), .D (nx8363), .CLK (clk), .R (rst)) ;
    mux21_ni ix8364 (.Y (nx8363), .A0 (camera_module_cache_ram_179__2), .A1 (
             nx35232), .S0 (nx34880)) ;
    dffr camera_module_cache_reg_ram_163__2 (.Q (camera_module_cache_ram_163__2)
         , .QB (\$dummy [600]), .D (nx8373), .CLK (clk), .R (rst)) ;
    mux21_ni ix8374 (.Y (nx8373), .A0 (camera_module_cache_ram_163__2), .A1 (
             nx35232), .S0 (nx34884)) ;
    aoi22 ix26743 (.Y (nx26742), .A0 (camera_module_cache_ram_195__2), .A1 (
          nx36298), .B0 (camera_module_cache_ram_211__2), .B1 (nx36338)) ;
    dffr camera_module_cache_reg_ram_195__2 (.Q (camera_module_cache_ram_195__2)
         , .QB (\$dummy [601]), .D (nx8353), .CLK (clk), .R (rst)) ;
    mux21_ni ix8354 (.Y (nx8353), .A0 (camera_module_cache_ram_195__2), .A1 (
             nx35232), .S0 (nx34876)) ;
    dffr camera_module_cache_reg_ram_211__2 (.Q (camera_module_cache_ram_211__2)
         , .QB (\$dummy [602]), .D (nx8343), .CLK (clk), .R (rst)) ;
    mux21_ni ix8344 (.Y (nx8343), .A0 (camera_module_cache_ram_211__2), .A1 (
             nx35232), .S0 (nx34872)) ;
    aoi22 ix26751 (.Y (nx26750), .A0 (camera_module_cache_ram_227__2), .A1 (
          nx36378), .B0 (camera_module_cache_ram_243__2), .B1 (nx36418)) ;
    dffr camera_module_cache_reg_ram_227__2 (.Q (camera_module_cache_ram_227__2)
         , .QB (\$dummy [603]), .D (nx8333), .CLK (clk), .R (rst)) ;
    mux21_ni ix8334 (.Y (nx8333), .A0 (camera_module_cache_ram_227__2), .A1 (
             nx35232), .S0 (nx34868)) ;
    dffr camera_module_cache_reg_ram_243__2 (.Q (camera_module_cache_ram_243__2)
         , .QB (\$dummy [604]), .D (nx8323), .CLK (clk), .R (rst)) ;
    mux21_ni ix8324 (.Y (nx8323), .A0 (camera_module_cache_ram_243__2), .A1 (
             nx35234), .S0 (nx34864)) ;
    nand04 ix10839 (.Y (nx10838), .A0 (nx26761), .A1 (nx26843), .A2 (nx26943), .A3 (
           nx27032)) ;
    oai21 ix26762 (.Y (nx26761), .A0 (nx10828), .A1 (nx10750), .B0 (nx36464)) ;
    nand04 ix10829 (.Y (nx10828), .A0 (nx26765), .A1 (nx26774), .A2 (nx26782), .A3 (
           nx26792)) ;
    aoi22 ix26766 (.Y (nx26765), .A0 (camera_module_cache_ram_4__2), .A1 (
          nx35818), .B0 (camera_module_cache_ram_20__2), .B1 (nx35858)) ;
    dffr camera_module_cache_reg_ram_4__2 (.Q (camera_module_cache_ram_4__2), .QB (
         \$dummy [605]), .D (nx8313), .CLK (clk), .R (rst)) ;
    mux21_ni ix8314 (.Y (nx8313), .A0 (camera_module_cache_ram_4__2), .A1 (
             nx35234), .S0 (nx34854)) ;
    dffr camera_module_cache_reg_ram_20__2 (.Q (camera_module_cache_ram_20__2), 
         .QB (\$dummy [606]), .D (nx8303), .CLK (clk), .R (rst)) ;
    mux21_ni ix8304 (.Y (nx8303), .A0 (camera_module_cache_ram_20__2), .A1 (
             nx35234), .S0 (nx34850)) ;
    aoi22 ix26775 (.Y (nx26774), .A0 (camera_module_cache_ram_36__2), .A1 (
          nx35898), .B0 (camera_module_cache_ram_52__2), .B1 (nx35938)) ;
    dffr camera_module_cache_reg_ram_36__2 (.Q (camera_module_cache_ram_36__2), 
         .QB (\$dummy [607]), .D (nx8293), .CLK (clk), .R (rst)) ;
    mux21_ni ix8294 (.Y (nx8293), .A0 (camera_module_cache_ram_36__2), .A1 (
             nx35234), .S0 (nx34846)) ;
    dffr camera_module_cache_reg_ram_52__2 (.Q (camera_module_cache_ram_52__2), 
         .QB (\$dummy [608]), .D (nx8283), .CLK (clk), .R (rst)) ;
    mux21_ni ix8284 (.Y (nx8283), .A0 (camera_module_cache_ram_52__2), .A1 (
             nx35234), .S0 (nx34842)) ;
    aoi22 ix26783 (.Y (nx26782), .A0 (camera_module_cache_ram_68__2), .A1 (
          nx35978), .B0 (camera_module_cache_ram_84__2), .B1 (nx36018)) ;
    dffr camera_module_cache_reg_ram_68__2 (.Q (camera_module_cache_ram_68__2), 
         .QB (\$dummy [609]), .D (nx8273), .CLK (clk), .R (rst)) ;
    mux21_ni ix8274 (.Y (nx8273), .A0 (camera_module_cache_ram_68__2), .A1 (
             nx35234), .S0 (nx34838)) ;
    dffr camera_module_cache_reg_ram_84__2 (.Q (camera_module_cache_ram_84__2), 
         .QB (\$dummy [610]), .D (nx8263), .CLK (clk), .R (rst)) ;
    mux21_ni ix8264 (.Y (nx8263), .A0 (camera_module_cache_ram_84__2), .A1 (
             nx35234), .S0 (nx34834)) ;
    aoi22 ix26793 (.Y (nx26792), .A0 (camera_module_cache_ram_116__2), .A1 (
          nx36058), .B0 (camera_module_cache_ram_100__2), .B1 (nx36098)) ;
    dffr camera_module_cache_reg_ram_116__2 (.Q (camera_module_cache_ram_116__2)
         , .QB (\$dummy [611]), .D (nx8243), .CLK (clk), .R (rst)) ;
    mux21_ni ix8244 (.Y (nx8243), .A0 (camera_module_cache_ram_116__2), .A1 (
             nx35236), .S0 (nx34826)) ;
    dffr camera_module_cache_reg_ram_100__2 (.Q (camera_module_cache_ram_100__2)
         , .QB (\$dummy [612]), .D (nx8253), .CLK (clk), .R (rst)) ;
    mux21_ni ix8254 (.Y (nx8253), .A0 (camera_module_cache_ram_100__2), .A1 (
             nx35236), .S0 (nx34830)) ;
    nand04 ix10751 (.Y (nx10750), .A0 (nx26803), .A1 (nx26813), .A2 (nx26822), .A3 (
           nx26831)) ;
    aoi22 ix26804 (.Y (nx26803), .A0 (camera_module_cache_ram_132__2), .A1 (
          nx36138), .B0 (camera_module_cache_ram_148__2), .B1 (nx36178)) ;
    dffr camera_module_cache_reg_ram_132__2 (.Q (camera_module_cache_ram_132__2)
         , .QB (\$dummy [613]), .D (nx8233), .CLK (clk), .R (rst)) ;
    mux21_ni ix8234 (.Y (nx8233), .A0 (camera_module_cache_ram_132__2), .A1 (
             nx35236), .S0 (nx34822)) ;
    dffr camera_module_cache_reg_ram_148__2 (.Q (camera_module_cache_ram_148__2)
         , .QB (\$dummy [614]), .D (nx8223), .CLK (clk), .R (rst)) ;
    mux21_ni ix8224 (.Y (nx8223), .A0 (camera_module_cache_ram_148__2), .A1 (
             nx35236), .S0 (nx34818)) ;
    aoi22 ix26814 (.Y (nx26813), .A0 (camera_module_cache_ram_180__2), .A1 (
          nx36218), .B0 (camera_module_cache_ram_164__2), .B1 (nx36258)) ;
    dffr camera_module_cache_reg_ram_180__2 (.Q (camera_module_cache_ram_180__2)
         , .QB (\$dummy [615]), .D (nx8203), .CLK (clk), .R (rst)) ;
    mux21_ni ix8204 (.Y (nx8203), .A0 (camera_module_cache_ram_180__2), .A1 (
             nx35236), .S0 (nx34810)) ;
    dffr camera_module_cache_reg_ram_164__2 (.Q (camera_module_cache_ram_164__2)
         , .QB (\$dummy [616]), .D (nx8213), .CLK (clk), .R (rst)) ;
    mux21_ni ix8214 (.Y (nx8213), .A0 (camera_module_cache_ram_164__2), .A1 (
             nx35236), .S0 (nx34814)) ;
    aoi22 ix26823 (.Y (nx26822), .A0 (camera_module_cache_ram_196__2), .A1 (
          nx36298), .B0 (camera_module_cache_ram_212__2), .B1 (nx36338)) ;
    dffr camera_module_cache_reg_ram_196__2 (.Q (camera_module_cache_ram_196__2)
         , .QB (\$dummy [617]), .D (nx8193), .CLK (clk), .R (rst)) ;
    mux21_ni ix8194 (.Y (nx8193), .A0 (camera_module_cache_ram_196__2), .A1 (
             nx35236), .S0 (nx34806)) ;
    dffr camera_module_cache_reg_ram_212__2 (.Q (camera_module_cache_ram_212__2)
         , .QB (\$dummy [618]), .D (nx8183), .CLK (clk), .R (rst)) ;
    mux21_ni ix8184 (.Y (nx8183), .A0 (camera_module_cache_ram_212__2), .A1 (
             nx35238), .S0 (nx34802)) ;
    aoi22 ix26832 (.Y (nx26831), .A0 (camera_module_cache_ram_228__2), .A1 (
          nx36378), .B0 (camera_module_cache_ram_244__2), .B1 (nx36418)) ;
    dffr camera_module_cache_reg_ram_228__2 (.Q (camera_module_cache_ram_228__2)
         , .QB (\$dummy [619]), .D (nx8173), .CLK (clk), .R (rst)) ;
    mux21_ni ix8174 (.Y (nx8173), .A0 (camera_module_cache_ram_228__2), .A1 (
             nx35238), .S0 (nx34798)) ;
    dffr camera_module_cache_reg_ram_244__2 (.Q (camera_module_cache_ram_244__2)
         , .QB (\$dummy [620]), .D (nx8163), .CLK (clk), .R (rst)) ;
    mux21_ni ix8164 (.Y (nx8163), .A0 (camera_module_cache_ram_244__2), .A1 (
             nx35238), .S0 (nx34794)) ;
    oai21 ix26844 (.Y (nx26843), .A0 (nx10666), .A1 (nx10588), .B0 (nx36468)) ;
    nand04 ix10667 (.Y (nx10666), .A0 (nx26847), .A1 (nx26859), .A2 (nx26871), .A3 (
           nx26883)) ;
    aoi22 ix26848 (.Y (nx26847), .A0 (camera_module_cache_ram_5__2), .A1 (
          nx35818), .B0 (camera_module_cache_ram_21__2), .B1 (nx35858)) ;
    dffr camera_module_cache_reg_ram_5__2 (.Q (camera_module_cache_ram_5__2), .QB (
         \$dummy [621]), .D (nx8153), .CLK (clk), .R (rst)) ;
    mux21_ni ix8154 (.Y (nx8153), .A0 (camera_module_cache_ram_5__2), .A1 (
             nx35238), .S0 (nx34784)) ;
    dffr camera_module_cache_reg_ram_21__2 (.Q (camera_module_cache_ram_21__2), 
         .QB (\$dummy [622]), .D (nx8143), .CLK (clk), .R (rst)) ;
    mux21_ni ix8144 (.Y (nx8143), .A0 (camera_module_cache_ram_21__2), .A1 (
             nx35238), .S0 (nx34780)) ;
    aoi22 ix26860 (.Y (nx26859), .A0 (camera_module_cache_ram_37__2), .A1 (
          nx35898), .B0 (camera_module_cache_ram_53__2), .B1 (nx35938)) ;
    dffr camera_module_cache_reg_ram_37__2 (.Q (camera_module_cache_ram_37__2), 
         .QB (\$dummy [623]), .D (nx8133), .CLK (clk), .R (rst)) ;
    mux21_ni ix8134 (.Y (nx8133), .A0 (camera_module_cache_ram_37__2), .A1 (
             nx35238), .S0 (nx34776)) ;
    dffr camera_module_cache_reg_ram_53__2 (.Q (camera_module_cache_ram_53__2), 
         .QB (\$dummy [624]), .D (nx8123), .CLK (clk), .R (rst)) ;
    mux21_ni ix8124 (.Y (nx8123), .A0 (camera_module_cache_ram_53__2), .A1 (
             nx35238), .S0 (nx34772)) ;
    aoi22 ix26872 (.Y (nx26871), .A0 (camera_module_cache_ram_69__2), .A1 (
          nx35978), .B0 (camera_module_cache_ram_85__2), .B1 (nx36018)) ;
    dffr camera_module_cache_reg_ram_69__2 (.Q (camera_module_cache_ram_69__2), 
         .QB (\$dummy [625]), .D (nx8113), .CLK (clk), .R (rst)) ;
    mux21_ni ix8114 (.Y (nx8113), .A0 (camera_module_cache_ram_69__2), .A1 (
             nx35240), .S0 (nx34768)) ;
    dffr camera_module_cache_reg_ram_85__2 (.Q (camera_module_cache_ram_85__2), 
         .QB (\$dummy [626]), .D (nx8103), .CLK (clk), .R (rst)) ;
    mux21_ni ix8104 (.Y (nx8103), .A0 (camera_module_cache_ram_85__2), .A1 (
             nx35240), .S0 (nx34764)) ;
    aoi22 ix26884 (.Y (nx26883), .A0 (camera_module_cache_ram_117__2), .A1 (
          nx36058), .B0 (camera_module_cache_ram_101__2), .B1 (nx36098)) ;
    dffr camera_module_cache_reg_ram_117__2 (.Q (camera_module_cache_ram_117__2)
         , .QB (\$dummy [627]), .D (nx8083), .CLK (clk), .R (rst)) ;
    mux21_ni ix8084 (.Y (nx8083), .A0 (camera_module_cache_ram_117__2), .A1 (
             nx35240), .S0 (nx34756)) ;
    dffr camera_module_cache_reg_ram_101__2 (.Q (camera_module_cache_ram_101__2)
         , .QB (\$dummy [628]), .D (nx8093), .CLK (clk), .R (rst)) ;
    mux21_ni ix8094 (.Y (nx8093), .A0 (camera_module_cache_ram_101__2), .A1 (
             nx35240), .S0 (nx34760)) ;
    nand04 ix10589 (.Y (nx10588), .A0 (nx26895), .A1 (nx26907), .A2 (nx26919), .A3 (
           nx26931)) ;
    aoi22 ix26896 (.Y (nx26895), .A0 (camera_module_cache_ram_133__2), .A1 (
          nx36138), .B0 (camera_module_cache_ram_149__2), .B1 (nx36178)) ;
    dffr camera_module_cache_reg_ram_133__2 (.Q (camera_module_cache_ram_133__2)
         , .QB (\$dummy [629]), .D (nx8073), .CLK (clk), .R (rst)) ;
    mux21_ni ix8074 (.Y (nx8073), .A0 (camera_module_cache_ram_133__2), .A1 (
             nx35240), .S0 (nx34752)) ;
    dffr camera_module_cache_reg_ram_149__2 (.Q (camera_module_cache_ram_149__2)
         , .QB (\$dummy [630]), .D (nx8063), .CLK (clk), .R (rst)) ;
    mux21_ni ix8064 (.Y (nx8063), .A0 (camera_module_cache_ram_149__2), .A1 (
             nx35240), .S0 (nx34748)) ;
    aoi22 ix26908 (.Y (nx26907), .A0 (camera_module_cache_ram_181__2), .A1 (
          nx36218), .B0 (camera_module_cache_ram_165__2), .B1 (nx36258)) ;
    dffr camera_module_cache_reg_ram_181__2 (.Q (camera_module_cache_ram_181__2)
         , .QB (\$dummy [631]), .D (nx8043), .CLK (clk), .R (rst)) ;
    mux21_ni ix8044 (.Y (nx8043), .A0 (camera_module_cache_ram_181__2), .A1 (
             nx35240), .S0 (nx34740)) ;
    dffr camera_module_cache_reg_ram_165__2 (.Q (camera_module_cache_ram_165__2)
         , .QB (\$dummy [632]), .D (nx8053), .CLK (clk), .R (rst)) ;
    mux21_ni ix8054 (.Y (nx8053), .A0 (camera_module_cache_ram_165__2), .A1 (
             nx35242), .S0 (nx34744)) ;
    aoi22 ix26920 (.Y (nx26919), .A0 (camera_module_cache_ram_197__2), .A1 (
          nx36298), .B0 (camera_module_cache_ram_213__2), .B1 (nx36338)) ;
    dffr camera_module_cache_reg_ram_197__2 (.Q (camera_module_cache_ram_197__2)
         , .QB (\$dummy [633]), .D (nx8033), .CLK (clk), .R (rst)) ;
    mux21_ni ix8034 (.Y (nx8033), .A0 (camera_module_cache_ram_197__2), .A1 (
             nx35242), .S0 (nx34736)) ;
    dffr camera_module_cache_reg_ram_213__2 (.Q (camera_module_cache_ram_213__2)
         , .QB (\$dummy [634]), .D (nx8023), .CLK (clk), .R (rst)) ;
    mux21_ni ix8024 (.Y (nx8023), .A0 (camera_module_cache_ram_213__2), .A1 (
             nx35242), .S0 (nx34732)) ;
    aoi22 ix26932 (.Y (nx26931), .A0 (camera_module_cache_ram_229__2), .A1 (
          nx36378), .B0 (camera_module_cache_ram_245__2), .B1 (nx36418)) ;
    dffr camera_module_cache_reg_ram_229__2 (.Q (camera_module_cache_ram_229__2)
         , .QB (\$dummy [635]), .D (nx8013), .CLK (clk), .R (rst)) ;
    mux21_ni ix8014 (.Y (nx8013), .A0 (camera_module_cache_ram_229__2), .A1 (
             nx35242), .S0 (nx34728)) ;
    dffr camera_module_cache_reg_ram_245__2 (.Q (camera_module_cache_ram_245__2)
         , .QB (\$dummy [636]), .D (nx8003), .CLK (clk), .R (rst)) ;
    mux21_ni ix8004 (.Y (nx8003), .A0 (camera_module_cache_ram_245__2), .A1 (
             nx35242), .S0 (nx34724)) ;
    oai21 ix26944 (.Y (nx26943), .A0 (nx10502), .A1 (nx10424), .B0 (nx36472)) ;
    nand04 ix10503 (.Y (nx10502), .A0 (nx26947), .A1 (nx26959), .A2 (nx26971), .A3 (
           nx26983)) ;
    aoi22 ix26948 (.Y (nx26947), .A0 (camera_module_cache_ram_6__2), .A1 (
          nx35820), .B0 (camera_module_cache_ram_22__2), .B1 (nx35860)) ;
    dffr camera_module_cache_reg_ram_6__2 (.Q (camera_module_cache_ram_6__2), .QB (
         \$dummy [637]), .D (nx7993), .CLK (clk), .R (rst)) ;
    mux21_ni ix7994 (.Y (nx7993), .A0 (camera_module_cache_ram_6__2), .A1 (
             nx35242), .S0 (nx34714)) ;
    dffr camera_module_cache_reg_ram_22__2 (.Q (camera_module_cache_ram_22__2), 
         .QB (\$dummy [638]), .D (nx7983), .CLK (clk), .R (rst)) ;
    mux21_ni ix7984 (.Y (nx7983), .A0 (camera_module_cache_ram_22__2), .A1 (
             nx35242), .S0 (nx34710)) ;
    aoi22 ix26960 (.Y (nx26959), .A0 (camera_module_cache_ram_38__2), .A1 (
          nx35900), .B0 (camera_module_cache_ram_54__2), .B1 (nx35940)) ;
    dffr camera_module_cache_reg_ram_38__2 (.Q (camera_module_cache_ram_38__2), 
         .QB (\$dummy [639]), .D (nx7973), .CLK (clk), .R (rst)) ;
    mux21_ni ix7974 (.Y (nx7973), .A0 (camera_module_cache_ram_38__2), .A1 (
             nx35244), .S0 (nx34706)) ;
    dffr camera_module_cache_reg_ram_54__2 (.Q (camera_module_cache_ram_54__2), 
         .QB (\$dummy [640]), .D (nx7963), .CLK (clk), .R (rst)) ;
    mux21_ni ix7964 (.Y (nx7963), .A0 (camera_module_cache_ram_54__2), .A1 (
             nx35244), .S0 (nx34702)) ;
    aoi22 ix26972 (.Y (nx26971), .A0 (camera_module_cache_ram_70__2), .A1 (
          nx35980), .B0 (camera_module_cache_ram_86__2), .B1 (nx36020)) ;
    dffr camera_module_cache_reg_ram_70__2 (.Q (camera_module_cache_ram_70__2), 
         .QB (\$dummy [641]), .D (nx7953), .CLK (clk), .R (rst)) ;
    mux21_ni ix7954 (.Y (nx7953), .A0 (camera_module_cache_ram_70__2), .A1 (
             nx35244), .S0 (nx34698)) ;
    dffr camera_module_cache_reg_ram_86__2 (.Q (camera_module_cache_ram_86__2), 
         .QB (\$dummy [642]), .D (nx7943), .CLK (clk), .R (rst)) ;
    mux21_ni ix7944 (.Y (nx7943), .A0 (camera_module_cache_ram_86__2), .A1 (
             nx35244), .S0 (nx34694)) ;
    aoi22 ix26984 (.Y (nx26983), .A0 (camera_module_cache_ram_118__2), .A1 (
          nx36060), .B0 (camera_module_cache_ram_102__2), .B1 (nx36100)) ;
    dffr camera_module_cache_reg_ram_118__2 (.Q (camera_module_cache_ram_118__2)
         , .QB (\$dummy [643]), .D (nx7923), .CLK (clk), .R (rst)) ;
    mux21_ni ix7924 (.Y (nx7923), .A0 (camera_module_cache_ram_118__2), .A1 (
             nx35244), .S0 (nx34686)) ;
    dffr camera_module_cache_reg_ram_102__2 (.Q (camera_module_cache_ram_102__2)
         , .QB (\$dummy [644]), .D (nx7933), .CLK (clk), .R (rst)) ;
    mux21_ni ix7934 (.Y (nx7933), .A0 (camera_module_cache_ram_102__2), .A1 (
             nx35244), .S0 (nx34690)) ;
    nand04 ix10425 (.Y (nx10424), .A0 (nx26993), .A1 (nx27004), .A2 (nx27013), .A3 (
           nx27023)) ;
    aoi22 ix26994 (.Y (nx26993), .A0 (camera_module_cache_ram_134__2), .A1 (
          nx36140), .B0 (camera_module_cache_ram_150__2), .B1 (nx36180)) ;
    dffr camera_module_cache_reg_ram_134__2 (.Q (camera_module_cache_ram_134__2)
         , .QB (\$dummy [645]), .D (nx7913), .CLK (clk), .R (rst)) ;
    mux21_ni ix7914 (.Y (nx7913), .A0 (camera_module_cache_ram_134__2), .A1 (
             nx35244), .S0 (nx34682)) ;
    dffr camera_module_cache_reg_ram_150__2 (.Q (camera_module_cache_ram_150__2)
         , .QB (\$dummy [646]), .D (nx7903), .CLK (clk), .R (rst)) ;
    mux21_ni ix7904 (.Y (nx7903), .A0 (camera_module_cache_ram_150__2), .A1 (
             nx35246), .S0 (nx34678)) ;
    aoi22 ix27005 (.Y (nx27004), .A0 (camera_module_cache_ram_182__2), .A1 (
          nx36220), .B0 (camera_module_cache_ram_166__2), .B1 (nx36260)) ;
    dffr camera_module_cache_reg_ram_182__2 (.Q (camera_module_cache_ram_182__2)
         , .QB (\$dummy [647]), .D (nx7883), .CLK (clk), .R (rst)) ;
    mux21_ni ix7884 (.Y (nx7883), .A0 (camera_module_cache_ram_182__2), .A1 (
             nx35246), .S0 (nx34670)) ;
    dffr camera_module_cache_reg_ram_166__2 (.Q (camera_module_cache_ram_166__2)
         , .QB (\$dummy [648]), .D (nx7893), .CLK (clk), .R (rst)) ;
    mux21_ni ix7894 (.Y (nx7893), .A0 (camera_module_cache_ram_166__2), .A1 (
             nx35246), .S0 (nx34674)) ;
    aoi22 ix27014 (.Y (nx27013), .A0 (camera_module_cache_ram_198__2), .A1 (
          nx36300), .B0 (camera_module_cache_ram_214__2), .B1 (nx36340)) ;
    dffr camera_module_cache_reg_ram_198__2 (.Q (camera_module_cache_ram_198__2)
         , .QB (\$dummy [649]), .D (nx7873), .CLK (clk), .R (rst)) ;
    mux21_ni ix7874 (.Y (nx7873), .A0 (camera_module_cache_ram_198__2), .A1 (
             nx35246), .S0 (nx34666)) ;
    dffr camera_module_cache_reg_ram_214__2 (.Q (camera_module_cache_ram_214__2)
         , .QB (\$dummy [650]), .D (nx7863), .CLK (clk), .R (rst)) ;
    mux21_ni ix7864 (.Y (nx7863), .A0 (camera_module_cache_ram_214__2), .A1 (
             nx35246), .S0 (nx34662)) ;
    aoi22 ix27024 (.Y (nx27023), .A0 (camera_module_cache_ram_230__2), .A1 (
          nx36380), .B0 (camera_module_cache_ram_246__2), .B1 (nx36420)) ;
    dffr camera_module_cache_reg_ram_230__2 (.Q (camera_module_cache_ram_230__2)
         , .QB (\$dummy [651]), .D (nx7853), .CLK (clk), .R (rst)) ;
    mux21_ni ix7854 (.Y (nx7853), .A0 (camera_module_cache_ram_230__2), .A1 (
             nx35246), .S0 (nx34658)) ;
    dffr camera_module_cache_reg_ram_246__2 (.Q (camera_module_cache_ram_246__2)
         , .QB (\$dummy [652]), .D (nx7843), .CLK (clk), .R (rst)) ;
    mux21_ni ix7844 (.Y (nx7843), .A0 (camera_module_cache_ram_246__2), .A1 (
             nx35246), .S0 (nx34654)) ;
    oai21 ix27033 (.Y (nx27032), .A0 (nx10340), .A1 (nx10262), .B0 (nx36476)) ;
    nand04 ix10341 (.Y (nx10340), .A0 (nx27035), .A1 (nx27045), .A2 (nx27054), .A3 (
           nx27065)) ;
    aoi22 ix27036 (.Y (nx27035), .A0 (camera_module_cache_ram_7__2), .A1 (
          nx35820), .B0 (camera_module_cache_ram_23__2), .B1 (nx35860)) ;
    dffr camera_module_cache_reg_ram_7__2 (.Q (camera_module_cache_ram_7__2), .QB (
         \$dummy [653]), .D (nx7833), .CLK (clk), .R (rst)) ;
    mux21_ni ix7834 (.Y (nx7833), .A0 (camera_module_cache_ram_7__2), .A1 (
             nx35248), .S0 (nx34644)) ;
    dffr camera_module_cache_reg_ram_23__2 (.Q (camera_module_cache_ram_23__2), 
         .QB (\$dummy [654]), .D (nx7823), .CLK (clk), .R (rst)) ;
    mux21_ni ix7824 (.Y (nx7823), .A0 (camera_module_cache_ram_23__2), .A1 (
             nx35248), .S0 (nx34640)) ;
    aoi22 ix27046 (.Y (nx27045), .A0 (camera_module_cache_ram_39__2), .A1 (
          nx35900), .B0 (camera_module_cache_ram_55__2), .B1 (nx35940)) ;
    dffr camera_module_cache_reg_ram_39__2 (.Q (camera_module_cache_ram_39__2), 
         .QB (\$dummy [655]), .D (nx7813), .CLK (clk), .R (rst)) ;
    mux21_ni ix7814 (.Y (nx7813), .A0 (camera_module_cache_ram_39__2), .A1 (
             nx35248), .S0 (nx34636)) ;
    dffr camera_module_cache_reg_ram_55__2 (.Q (camera_module_cache_ram_55__2), 
         .QB (\$dummy [656]), .D (nx7803), .CLK (clk), .R (rst)) ;
    mux21_ni ix7804 (.Y (nx7803), .A0 (camera_module_cache_ram_55__2), .A1 (
             nx35248), .S0 (nx34632)) ;
    aoi22 ix27055 (.Y (nx27054), .A0 (camera_module_cache_ram_71__2), .A1 (
          nx35980), .B0 (camera_module_cache_ram_87__2), .B1 (nx36020)) ;
    dffr camera_module_cache_reg_ram_71__2 (.Q (camera_module_cache_ram_71__2), 
         .QB (\$dummy [657]), .D (nx7793), .CLK (clk), .R (rst)) ;
    mux21_ni ix7794 (.Y (nx7793), .A0 (camera_module_cache_ram_71__2), .A1 (
             nx35248), .S0 (nx34628)) ;
    dffr camera_module_cache_reg_ram_87__2 (.Q (camera_module_cache_ram_87__2), 
         .QB (\$dummy [658]), .D (nx7783), .CLK (clk), .R (rst)) ;
    mux21_ni ix7784 (.Y (nx7783), .A0 (camera_module_cache_ram_87__2), .A1 (
             nx35248), .S0 (nx34624)) ;
    aoi22 ix27066 (.Y (nx27065), .A0 (camera_module_cache_ram_119__2), .A1 (
          nx36060), .B0 (camera_module_cache_ram_103__2), .B1 (nx36100)) ;
    dffr camera_module_cache_reg_ram_119__2 (.Q (camera_module_cache_ram_119__2)
         , .QB (\$dummy [659]), .D (nx7763), .CLK (clk), .R (rst)) ;
    mux21_ni ix7764 (.Y (nx7763), .A0 (camera_module_cache_ram_119__2), .A1 (
             nx35248), .S0 (nx34616)) ;
    dffr camera_module_cache_reg_ram_103__2 (.Q (camera_module_cache_ram_103__2)
         , .QB (\$dummy [660]), .D (nx7773), .CLK (clk), .R (rst)) ;
    mux21_ni ix7774 (.Y (nx7773), .A0 (camera_module_cache_ram_103__2), .A1 (
             nx35250), .S0 (nx34620)) ;
    nand04 ix10263 (.Y (nx10262), .A0 (nx27076), .A1 (nx27088), .A2 (nx27097), .A3 (
           nx27105)) ;
    aoi22 ix27078 (.Y (nx27076), .A0 (camera_module_cache_ram_135__2), .A1 (
          nx36140), .B0 (camera_module_cache_ram_151__2), .B1 (nx36180)) ;
    dffr camera_module_cache_reg_ram_135__2 (.Q (camera_module_cache_ram_135__2)
         , .QB (\$dummy [661]), .D (nx7753), .CLK (clk), .R (rst)) ;
    mux21_ni ix7754 (.Y (nx7753), .A0 (camera_module_cache_ram_135__2), .A1 (
             nx35250), .S0 (nx34612)) ;
    dffr camera_module_cache_reg_ram_151__2 (.Q (camera_module_cache_ram_151__2)
         , .QB (\$dummy [662]), .D (nx7743), .CLK (clk), .R (rst)) ;
    mux21_ni ix7744 (.Y (nx7743), .A0 (camera_module_cache_ram_151__2), .A1 (
             nx35250), .S0 (nx34608)) ;
    aoi22 ix27089 (.Y (nx27088), .A0 (camera_module_cache_ram_183__2), .A1 (
          nx36220), .B0 (camera_module_cache_ram_167__2), .B1 (nx36260)) ;
    dffr camera_module_cache_reg_ram_183__2 (.Q (camera_module_cache_ram_183__2)
         , .QB (\$dummy [663]), .D (nx7723), .CLK (clk), .R (rst)) ;
    mux21_ni ix7724 (.Y (nx7723), .A0 (camera_module_cache_ram_183__2), .A1 (
             nx35250), .S0 (nx34600)) ;
    dffr camera_module_cache_reg_ram_167__2 (.Q (camera_module_cache_ram_167__2)
         , .QB (\$dummy [664]), .D (nx7733), .CLK (clk), .R (rst)) ;
    mux21_ni ix7734 (.Y (nx7733), .A0 (camera_module_cache_ram_167__2), .A1 (
             nx35250), .S0 (nx34604)) ;
    aoi22 ix27098 (.Y (nx27097), .A0 (camera_module_cache_ram_199__2), .A1 (
          nx36300), .B0 (camera_module_cache_ram_215__2), .B1 (nx36340)) ;
    dffr camera_module_cache_reg_ram_199__2 (.Q (camera_module_cache_ram_199__2)
         , .QB (\$dummy [665]), .D (nx7713), .CLK (clk), .R (rst)) ;
    mux21_ni ix7714 (.Y (nx7713), .A0 (camera_module_cache_ram_199__2), .A1 (
             nx35250), .S0 (nx34596)) ;
    dffr camera_module_cache_reg_ram_215__2 (.Q (camera_module_cache_ram_215__2)
         , .QB (\$dummy [666]), .D (nx7703), .CLK (clk), .R (rst)) ;
    mux21_ni ix7704 (.Y (nx7703), .A0 (camera_module_cache_ram_215__2), .A1 (
             nx35250), .S0 (nx34592)) ;
    aoi22 ix27106 (.Y (nx27105), .A0 (camera_module_cache_ram_231__2), .A1 (
          nx36380), .B0 (camera_module_cache_ram_247__2), .B1 (nx36420)) ;
    dffr camera_module_cache_reg_ram_231__2 (.Q (camera_module_cache_ram_231__2)
         , .QB (\$dummy [667]), .D (nx7693), .CLK (clk), .R (rst)) ;
    mux21_ni ix7694 (.Y (nx7693), .A0 (camera_module_cache_ram_231__2), .A1 (
             nx35252), .S0 (nx34588)) ;
    dffr camera_module_cache_reg_ram_247__2 (.Q (camera_module_cache_ram_247__2)
         , .QB (\$dummy [668]), .D (nx7683), .CLK (clk), .R (rst)) ;
    mux21_ni ix7684 (.Y (nx7683), .A0 (camera_module_cache_ram_247__2), .A1 (
             nx35252), .S0 (nx34584)) ;
    nand04 ix10183 (.Y (nx10182), .A0 (nx27115), .A1 (nx27197), .A2 (nx27265), .A3 (
           nx27333)) ;
    oai21 ix27116 (.Y (nx27115), .A0 (nx10172), .A1 (nx10094), .B0 (nx36480)) ;
    nand04 ix10173 (.Y (nx10172), .A0 (nx27119), .A1 (nx27131), .A2 (nx27142), .A3 (
           nx27152)) ;
    aoi22 ix27120 (.Y (nx27119), .A0 (camera_module_cache_ram_8__2), .A1 (
          nx35820), .B0 (camera_module_cache_ram_24__2), .B1 (nx35860)) ;
    dffr camera_module_cache_reg_ram_8__2 (.Q (camera_module_cache_ram_8__2), .QB (
         \$dummy [669]), .D (nx7673), .CLK (clk), .R (rst)) ;
    mux21_ni ix7674 (.Y (nx7673), .A0 (camera_module_cache_ram_8__2), .A1 (
             nx35252), .S0 (nx34574)) ;
    dffr camera_module_cache_reg_ram_24__2 (.Q (camera_module_cache_ram_24__2), 
         .QB (\$dummy [670]), .D (nx7663), .CLK (clk), .R (rst)) ;
    mux21_ni ix7664 (.Y (nx7663), .A0 (camera_module_cache_ram_24__2), .A1 (
             nx35252), .S0 (nx34570)) ;
    aoi22 ix27132 (.Y (nx27131), .A0 (camera_module_cache_ram_40__2), .A1 (
          nx35900), .B0 (camera_module_cache_ram_56__2), .B1 (nx35940)) ;
    dffr camera_module_cache_reg_ram_40__2 (.Q (camera_module_cache_ram_40__2), 
         .QB (\$dummy [671]), .D (nx7653), .CLK (clk), .R (rst)) ;
    mux21_ni ix7654 (.Y (nx7653), .A0 (camera_module_cache_ram_40__2), .A1 (
             nx35252), .S0 (nx34566)) ;
    dffr camera_module_cache_reg_ram_56__2 (.Q (camera_module_cache_ram_56__2), 
         .QB (\$dummy [672]), .D (nx7643), .CLK (clk), .R (rst)) ;
    mux21_ni ix7644 (.Y (nx7643), .A0 (camera_module_cache_ram_56__2), .A1 (
             nx35252), .S0 (nx34562)) ;
    aoi22 ix27144 (.Y (nx27142), .A0 (camera_module_cache_ram_72__2), .A1 (
          nx35980), .B0 (camera_module_cache_ram_88__2), .B1 (nx36020)) ;
    dffr camera_module_cache_reg_ram_72__2 (.Q (camera_module_cache_ram_72__2), 
         .QB (\$dummy [673]), .D (nx7633), .CLK (clk), .R (rst)) ;
    mux21_ni ix7634 (.Y (nx7633), .A0 (camera_module_cache_ram_72__2), .A1 (
             nx35252), .S0 (nx34558)) ;
    dffr camera_module_cache_reg_ram_88__2 (.Q (camera_module_cache_ram_88__2), 
         .QB (\$dummy [674]), .D (nx7623), .CLK (clk), .R (rst)) ;
    mux21_ni ix7624 (.Y (nx7623), .A0 (camera_module_cache_ram_88__2), .A1 (
             nx35254), .S0 (nx34554)) ;
    aoi22 ix27153 (.Y (nx27152), .A0 (camera_module_cache_ram_120__2), .A1 (
          nx36060), .B0 (camera_module_cache_ram_104__2), .B1 (nx36100)) ;
    dffr camera_module_cache_reg_ram_120__2 (.Q (camera_module_cache_ram_120__2)
         , .QB (\$dummy [675]), .D (nx7603), .CLK (clk), .R (rst)) ;
    mux21_ni ix7604 (.Y (nx7603), .A0 (camera_module_cache_ram_120__2), .A1 (
             nx35254), .S0 (nx34546)) ;
    dffr camera_module_cache_reg_ram_104__2 (.Q (camera_module_cache_ram_104__2)
         , .QB (\$dummy [676]), .D (nx7613), .CLK (clk), .R (rst)) ;
    mux21_ni ix7614 (.Y (nx7613), .A0 (camera_module_cache_ram_104__2), .A1 (
             nx35254), .S0 (nx34550)) ;
    nand04 ix10095 (.Y (nx10094), .A0 (nx27163), .A1 (nx27173), .A2 (nx27181), .A3 (
           nx27189)) ;
    aoi22 ix27164 (.Y (nx27163), .A0 (camera_module_cache_ram_136__2), .A1 (
          nx36140), .B0 (camera_module_cache_ram_152__2), .B1 (nx36180)) ;
    dffr camera_module_cache_reg_ram_136__2 (.Q (camera_module_cache_ram_136__2)
         , .QB (\$dummy [677]), .D (nx7593), .CLK (clk), .R (rst)) ;
    mux21_ni ix7594 (.Y (nx7593), .A0 (camera_module_cache_ram_136__2), .A1 (
             nx35254), .S0 (nx34542)) ;
    dffr camera_module_cache_reg_ram_152__2 (.Q (camera_module_cache_ram_152__2)
         , .QB (\$dummy [678]), .D (nx7583), .CLK (clk), .R (rst)) ;
    mux21_ni ix7584 (.Y (nx7583), .A0 (camera_module_cache_ram_152__2), .A1 (
             nx35254), .S0 (nx34538)) ;
    aoi22 ix27174 (.Y (nx27173), .A0 (camera_module_cache_ram_184__2), .A1 (
          nx36220), .B0 (camera_module_cache_ram_168__2), .B1 (nx36260)) ;
    dffr camera_module_cache_reg_ram_184__2 (.Q (camera_module_cache_ram_184__2)
         , .QB (\$dummy [679]), .D (nx7563), .CLK (clk), .R (rst)) ;
    mux21_ni ix7564 (.Y (nx7563), .A0 (camera_module_cache_ram_184__2), .A1 (
             nx35254), .S0 (nx34530)) ;
    dffr camera_module_cache_reg_ram_168__2 (.Q (camera_module_cache_ram_168__2)
         , .QB (\$dummy [680]), .D (nx7573), .CLK (clk), .R (rst)) ;
    mux21_ni ix7574 (.Y (nx7573), .A0 (camera_module_cache_ram_168__2), .A1 (
             nx35254), .S0 (nx34534)) ;
    aoi22 ix27182 (.Y (nx27181), .A0 (camera_module_cache_ram_200__2), .A1 (
          nx36300), .B0 (camera_module_cache_ram_216__2), .B1 (nx36340)) ;
    dffr camera_module_cache_reg_ram_200__2 (.Q (camera_module_cache_ram_200__2)
         , .QB (\$dummy [681]), .D (nx7553), .CLK (clk), .R (rst)) ;
    mux21_ni ix7554 (.Y (nx7553), .A0 (camera_module_cache_ram_200__2), .A1 (
             nx35256), .S0 (nx34526)) ;
    dffr camera_module_cache_reg_ram_216__2 (.Q (camera_module_cache_ram_216__2)
         , .QB (\$dummy [682]), .D (nx7543), .CLK (clk), .R (rst)) ;
    mux21_ni ix7544 (.Y (nx7543), .A0 (camera_module_cache_ram_216__2), .A1 (
             nx35256), .S0 (nx34522)) ;
    aoi22 ix27190 (.Y (nx27189), .A0 (camera_module_cache_ram_232__2), .A1 (
          nx36380), .B0 (camera_module_cache_ram_248__2), .B1 (nx36420)) ;
    dffr camera_module_cache_reg_ram_232__2 (.Q (camera_module_cache_ram_232__2)
         , .QB (\$dummy [683]), .D (nx7533), .CLK (clk), .R (rst)) ;
    mux21_ni ix7534 (.Y (nx7533), .A0 (camera_module_cache_ram_232__2), .A1 (
             nx35256), .S0 (nx34518)) ;
    dffr camera_module_cache_reg_ram_248__2 (.Q (camera_module_cache_ram_248__2)
         , .QB (\$dummy [684]), .D (nx7523), .CLK (clk), .R (rst)) ;
    mux21_ni ix7524 (.Y (nx7523), .A0 (camera_module_cache_ram_248__2), .A1 (
             nx35256), .S0 (nx34514)) ;
    oai21 ix27198 (.Y (nx27197), .A0 (nx10010), .A1 (nx9932), .B0 (nx36484)) ;
    nand04 ix10011 (.Y (nx10010), .A0 (nx27200), .A1 (nx27208), .A2 (nx27216), .A3 (
           nx27224)) ;
    aoi22 ix27201 (.Y (nx27200), .A0 (camera_module_cache_ram_9__2), .A1 (
          nx35820), .B0 (camera_module_cache_ram_25__2), .B1 (nx35860)) ;
    dffr camera_module_cache_reg_ram_9__2 (.Q (camera_module_cache_ram_9__2), .QB (
         \$dummy [685]), .D (nx7513), .CLK (clk), .R (rst)) ;
    mux21_ni ix7514 (.Y (nx7513), .A0 (camera_module_cache_ram_9__2), .A1 (
             nx35256), .S0 (nx34504)) ;
    dffr camera_module_cache_reg_ram_25__2 (.Q (camera_module_cache_ram_25__2), 
         .QB (\$dummy [686]), .D (nx7503), .CLK (clk), .R (rst)) ;
    mux21_ni ix7504 (.Y (nx7503), .A0 (camera_module_cache_ram_25__2), .A1 (
             nx35256), .S0 (nx34500)) ;
    aoi22 ix27209 (.Y (nx27208), .A0 (camera_module_cache_ram_41__2), .A1 (
          nx35900), .B0 (camera_module_cache_ram_57__2), .B1 (nx35940)) ;
    dffr camera_module_cache_reg_ram_41__2 (.Q (camera_module_cache_ram_41__2), 
         .QB (\$dummy [687]), .D (nx7493), .CLK (clk), .R (rst)) ;
    mux21_ni ix7494 (.Y (nx7493), .A0 (camera_module_cache_ram_41__2), .A1 (
             nx35256), .S0 (nx34496)) ;
    dffr camera_module_cache_reg_ram_57__2 (.Q (camera_module_cache_ram_57__2), 
         .QB (\$dummy [688]), .D (nx7483), .CLK (clk), .R (rst)) ;
    mux21_ni ix7484 (.Y (nx7483), .A0 (camera_module_cache_ram_57__2), .A1 (
             nx35258), .S0 (nx34492)) ;
    aoi22 ix27217 (.Y (nx27216), .A0 (camera_module_cache_ram_73__2), .A1 (
          nx35980), .B0 (camera_module_cache_ram_89__2), .B1 (nx36020)) ;
    dffr camera_module_cache_reg_ram_73__2 (.Q (camera_module_cache_ram_73__2), 
         .QB (\$dummy [689]), .D (nx7473), .CLK (clk), .R (rst)) ;
    mux21_ni ix7474 (.Y (nx7473), .A0 (camera_module_cache_ram_73__2), .A1 (
             nx35258), .S0 (nx34488)) ;
    dffr camera_module_cache_reg_ram_89__2 (.Q (camera_module_cache_ram_89__2), 
         .QB (\$dummy [690]), .D (nx7463), .CLK (clk), .R (rst)) ;
    mux21_ni ix7464 (.Y (nx7463), .A0 (camera_module_cache_ram_89__2), .A1 (
             nx35258), .S0 (nx34484)) ;
    aoi22 ix27225 (.Y (nx27224), .A0 (camera_module_cache_ram_121__2), .A1 (
          nx36060), .B0 (camera_module_cache_ram_105__2), .B1 (nx36100)) ;
    dffr camera_module_cache_reg_ram_121__2 (.Q (camera_module_cache_ram_121__2)
         , .QB (\$dummy [691]), .D (nx7443), .CLK (clk), .R (rst)) ;
    mux21_ni ix7444 (.Y (nx7443), .A0 (camera_module_cache_ram_121__2), .A1 (
             nx35258), .S0 (nx34476)) ;
    dffr camera_module_cache_reg_ram_105__2 (.Q (camera_module_cache_ram_105__2)
         , .QB (\$dummy [692]), .D (nx7453), .CLK (clk), .R (rst)) ;
    mux21_ni ix7454 (.Y (nx7453), .A0 (camera_module_cache_ram_105__2), .A1 (
             nx35258), .S0 (nx34480)) ;
    nand04 ix9933 (.Y (nx9932), .A0 (nx27233), .A1 (nx27241), .A2 (nx27249), .A3 (
           nx27257)) ;
    aoi22 ix27234 (.Y (nx27233), .A0 (camera_module_cache_ram_137__2), .A1 (
          nx36140), .B0 (camera_module_cache_ram_153__2), .B1 (nx36180)) ;
    dffr camera_module_cache_reg_ram_137__2 (.Q (camera_module_cache_ram_137__2)
         , .QB (\$dummy [693]), .D (nx7433), .CLK (clk), .R (rst)) ;
    mux21_ni ix7434 (.Y (nx7433), .A0 (camera_module_cache_ram_137__2), .A1 (
             nx35258), .S0 (nx34472)) ;
    dffr camera_module_cache_reg_ram_153__2 (.Q (camera_module_cache_ram_153__2)
         , .QB (\$dummy [694]), .D (nx7423), .CLK (clk), .R (rst)) ;
    mux21_ni ix7424 (.Y (nx7423), .A0 (camera_module_cache_ram_153__2), .A1 (
             nx35258), .S0 (nx34468)) ;
    aoi22 ix27242 (.Y (nx27241), .A0 (camera_module_cache_ram_185__2), .A1 (
          nx36220), .B0 (camera_module_cache_ram_169__2), .B1 (nx36260)) ;
    dffr camera_module_cache_reg_ram_185__2 (.Q (camera_module_cache_ram_185__2)
         , .QB (\$dummy [695]), .D (nx7403), .CLK (clk), .R (rst)) ;
    mux21_ni ix7404 (.Y (nx7403), .A0 (camera_module_cache_ram_185__2), .A1 (
             nx35260), .S0 (nx34460)) ;
    dffr camera_module_cache_reg_ram_169__2 (.Q (camera_module_cache_ram_169__2)
         , .QB (\$dummy [696]), .D (nx7413), .CLK (clk), .R (rst)) ;
    mux21_ni ix7414 (.Y (nx7413), .A0 (camera_module_cache_ram_169__2), .A1 (
             nx35260), .S0 (nx34464)) ;
    aoi22 ix27250 (.Y (nx27249), .A0 (camera_module_cache_ram_201__2), .A1 (
          nx36300), .B0 (camera_module_cache_ram_217__2), .B1 (nx36340)) ;
    dffr camera_module_cache_reg_ram_201__2 (.Q (camera_module_cache_ram_201__2)
         , .QB (\$dummy [697]), .D (nx7393), .CLK (clk), .R (rst)) ;
    mux21_ni ix7394 (.Y (nx7393), .A0 (camera_module_cache_ram_201__2), .A1 (
             nx35260), .S0 (nx34456)) ;
    dffr camera_module_cache_reg_ram_217__2 (.Q (camera_module_cache_ram_217__2)
         , .QB (\$dummy [698]), .D (nx7383), .CLK (clk), .R (rst)) ;
    mux21_ni ix7384 (.Y (nx7383), .A0 (camera_module_cache_ram_217__2), .A1 (
             nx35260), .S0 (nx34452)) ;
    aoi22 ix27258 (.Y (nx27257), .A0 (camera_module_cache_ram_233__2), .A1 (
          nx36380), .B0 (camera_module_cache_ram_249__2), .B1 (nx36420)) ;
    dffr camera_module_cache_reg_ram_233__2 (.Q (camera_module_cache_ram_233__2)
         , .QB (\$dummy [699]), .D (nx7373), .CLK (clk), .R (rst)) ;
    mux21_ni ix7374 (.Y (nx7373), .A0 (camera_module_cache_ram_233__2), .A1 (
             nx35260), .S0 (nx34448)) ;
    dffr camera_module_cache_reg_ram_249__2 (.Q (camera_module_cache_ram_249__2)
         , .QB (\$dummy [700]), .D (nx7363), .CLK (clk), .R (rst)) ;
    mux21_ni ix7364 (.Y (nx7363), .A0 (camera_module_cache_ram_249__2), .A1 (
             nx35260), .S0 (nx34444)) ;
    oai21 ix27266 (.Y (nx27265), .A0 (nx9846), .A1 (nx9768), .B0 (nx36488)) ;
    nand04 ix9847 (.Y (nx9846), .A0 (nx27268), .A1 (nx27276), .A2 (nx27284), .A3 (
           nx27292)) ;
    aoi22 ix27269 (.Y (nx27268), .A0 (camera_module_cache_ram_10__2), .A1 (
          nx35820), .B0 (camera_module_cache_ram_26__2), .B1 (nx35860)) ;
    dffr camera_module_cache_reg_ram_10__2 (.Q (camera_module_cache_ram_10__2), 
         .QB (\$dummy [701]), .D (nx7353), .CLK (clk), .R (rst)) ;
    mux21_ni ix7354 (.Y (nx7353), .A0 (camera_module_cache_ram_10__2), .A1 (
             nx35260), .S0 (nx34434)) ;
    dffr camera_module_cache_reg_ram_26__2 (.Q (camera_module_cache_ram_26__2), 
         .QB (\$dummy [702]), .D (nx7343), .CLK (clk), .R (rst)) ;
    mux21_ni ix7344 (.Y (nx7343), .A0 (camera_module_cache_ram_26__2), .A1 (
             nx35262), .S0 (nx34430)) ;
    aoi22 ix27277 (.Y (nx27276), .A0 (camera_module_cache_ram_42__2), .A1 (
          nx35900), .B0 (camera_module_cache_ram_58__2), .B1 (nx35940)) ;
    dffr camera_module_cache_reg_ram_42__2 (.Q (camera_module_cache_ram_42__2), 
         .QB (\$dummy [703]), .D (nx7333), .CLK (clk), .R (rst)) ;
    mux21_ni ix7334 (.Y (nx7333), .A0 (camera_module_cache_ram_42__2), .A1 (
             nx35262), .S0 (nx34426)) ;
    dffr camera_module_cache_reg_ram_58__2 (.Q (camera_module_cache_ram_58__2), 
         .QB (\$dummy [704]), .D (nx7323), .CLK (clk), .R (rst)) ;
    mux21_ni ix7324 (.Y (nx7323), .A0 (camera_module_cache_ram_58__2), .A1 (
             nx35262), .S0 (nx34422)) ;
    aoi22 ix27285 (.Y (nx27284), .A0 (camera_module_cache_ram_74__2), .A1 (
          nx35980), .B0 (camera_module_cache_ram_90__2), .B1 (nx36020)) ;
    dffr camera_module_cache_reg_ram_74__2 (.Q (camera_module_cache_ram_74__2), 
         .QB (\$dummy [705]), .D (nx7313), .CLK (clk), .R (rst)) ;
    mux21_ni ix7314 (.Y (nx7313), .A0 (camera_module_cache_ram_74__2), .A1 (
             nx35262), .S0 (nx34418)) ;
    dffr camera_module_cache_reg_ram_90__2 (.Q (camera_module_cache_ram_90__2), 
         .QB (\$dummy [706]), .D (nx7303), .CLK (clk), .R (rst)) ;
    mux21_ni ix7304 (.Y (nx7303), .A0 (camera_module_cache_ram_90__2), .A1 (
             nx35262), .S0 (nx34414)) ;
    aoi22 ix27293 (.Y (nx27292), .A0 (camera_module_cache_ram_122__2), .A1 (
          nx36060), .B0 (camera_module_cache_ram_106__2), .B1 (nx36100)) ;
    dffr camera_module_cache_reg_ram_122__2 (.Q (camera_module_cache_ram_122__2)
         , .QB (\$dummy [707]), .D (nx7283), .CLK (clk), .R (rst)) ;
    mux21_ni ix7284 (.Y (nx7283), .A0 (camera_module_cache_ram_122__2), .A1 (
             nx35262), .S0 (nx34406)) ;
    dffr camera_module_cache_reg_ram_106__2 (.Q (camera_module_cache_ram_106__2)
         , .QB (\$dummy [708]), .D (nx7293), .CLK (clk), .R (rst)) ;
    mux21_ni ix7294 (.Y (nx7293), .A0 (camera_module_cache_ram_106__2), .A1 (
             nx35262), .S0 (nx34410)) ;
    nand04 ix9769 (.Y (nx9768), .A0 (nx27301), .A1 (nx27309), .A2 (nx27317), .A3 (
           nx27325)) ;
    aoi22 ix27302 (.Y (nx27301), .A0 (camera_module_cache_ram_138__2), .A1 (
          nx36140), .B0 (camera_module_cache_ram_154__2), .B1 (nx36180)) ;
    dffr camera_module_cache_reg_ram_138__2 (.Q (camera_module_cache_ram_138__2)
         , .QB (\$dummy [709]), .D (nx7273), .CLK (clk), .R (rst)) ;
    mux21_ni ix7274 (.Y (nx7273), .A0 (camera_module_cache_ram_138__2), .A1 (
             nx35264), .S0 (nx34402)) ;
    dffr camera_module_cache_reg_ram_154__2 (.Q (camera_module_cache_ram_154__2)
         , .QB (\$dummy [710]), .D (nx7263), .CLK (clk), .R (rst)) ;
    mux21_ni ix7264 (.Y (nx7263), .A0 (camera_module_cache_ram_154__2), .A1 (
             nx35264), .S0 (nx34398)) ;
    aoi22 ix27310 (.Y (nx27309), .A0 (camera_module_cache_ram_186__2), .A1 (
          nx36220), .B0 (camera_module_cache_ram_170__2), .B1 (nx36260)) ;
    dffr camera_module_cache_reg_ram_186__2 (.Q (camera_module_cache_ram_186__2)
         , .QB (\$dummy [711]), .D (nx7243), .CLK (clk), .R (rst)) ;
    mux21_ni ix7244 (.Y (nx7243), .A0 (camera_module_cache_ram_186__2), .A1 (
             nx35264), .S0 (nx34390)) ;
    dffr camera_module_cache_reg_ram_170__2 (.Q (camera_module_cache_ram_170__2)
         , .QB (\$dummy [712]), .D (nx7253), .CLK (clk), .R (rst)) ;
    mux21_ni ix7254 (.Y (nx7253), .A0 (camera_module_cache_ram_170__2), .A1 (
             nx35264), .S0 (nx34394)) ;
    aoi22 ix27318 (.Y (nx27317), .A0 (camera_module_cache_ram_202__2), .A1 (
          nx36300), .B0 (camera_module_cache_ram_218__2), .B1 (nx36340)) ;
    dffr camera_module_cache_reg_ram_202__2 (.Q (camera_module_cache_ram_202__2)
         , .QB (\$dummy [713]), .D (nx7233), .CLK (clk), .R (rst)) ;
    mux21_ni ix7234 (.Y (nx7233), .A0 (camera_module_cache_ram_202__2), .A1 (
             nx35264), .S0 (nx34386)) ;
    dffr camera_module_cache_reg_ram_218__2 (.Q (camera_module_cache_ram_218__2)
         , .QB (\$dummy [714]), .D (nx7223), .CLK (clk), .R (rst)) ;
    mux21_ni ix7224 (.Y (nx7223), .A0 (camera_module_cache_ram_218__2), .A1 (
             nx35264), .S0 (nx34382)) ;
    aoi22 ix27326 (.Y (nx27325), .A0 (camera_module_cache_ram_234__2), .A1 (
          nx36380), .B0 (camera_module_cache_ram_250__2), .B1 (nx36420)) ;
    dffr camera_module_cache_reg_ram_234__2 (.Q (camera_module_cache_ram_234__2)
         , .QB (\$dummy [715]), .D (nx7213), .CLK (clk), .R (rst)) ;
    mux21_ni ix7214 (.Y (nx7213), .A0 (camera_module_cache_ram_234__2), .A1 (
             nx35264), .S0 (nx34378)) ;
    dffr camera_module_cache_reg_ram_250__2 (.Q (camera_module_cache_ram_250__2)
         , .QB (\$dummy [716]), .D (nx7203), .CLK (clk), .R (rst)) ;
    mux21_ni ix7204 (.Y (nx7203), .A0 (camera_module_cache_ram_250__2), .A1 (
             nx35266), .S0 (nx34374)) ;
    oai21 ix27334 (.Y (nx27333), .A0 (nx9684), .A1 (nx9606), .B0 (nx36492)) ;
    nand04 ix9685 (.Y (nx9684), .A0 (nx27336), .A1 (nx27344), .A2 (nx27352), .A3 (
           nx27360)) ;
    aoi22 ix27337 (.Y (nx27336), .A0 (camera_module_cache_ram_11__2), .A1 (
          nx35820), .B0 (camera_module_cache_ram_27__2), .B1 (nx35860)) ;
    dffr camera_module_cache_reg_ram_11__2 (.Q (camera_module_cache_ram_11__2), 
         .QB (\$dummy [717]), .D (nx7193), .CLK (clk), .R (rst)) ;
    mux21_ni ix7194 (.Y (nx7193), .A0 (camera_module_cache_ram_11__2), .A1 (
             nx35266), .S0 (nx34364)) ;
    dffr camera_module_cache_reg_ram_27__2 (.Q (camera_module_cache_ram_27__2), 
         .QB (\$dummy [718]), .D (nx7183), .CLK (clk), .R (rst)) ;
    mux21_ni ix7184 (.Y (nx7183), .A0 (camera_module_cache_ram_27__2), .A1 (
             nx35266), .S0 (nx34360)) ;
    aoi22 ix27345 (.Y (nx27344), .A0 (camera_module_cache_ram_43__2), .A1 (
          nx35900), .B0 (camera_module_cache_ram_59__2), .B1 (nx35940)) ;
    dffr camera_module_cache_reg_ram_43__2 (.Q (camera_module_cache_ram_43__2), 
         .QB (\$dummy [719]), .D (nx7173), .CLK (clk), .R (rst)) ;
    mux21_ni ix7174 (.Y (nx7173), .A0 (camera_module_cache_ram_43__2), .A1 (
             nx35266), .S0 (nx34356)) ;
    dffr camera_module_cache_reg_ram_59__2 (.Q (camera_module_cache_ram_59__2), 
         .QB (\$dummy [720]), .D (nx7163), .CLK (clk), .R (rst)) ;
    mux21_ni ix7164 (.Y (nx7163), .A0 (camera_module_cache_ram_59__2), .A1 (
             nx35266), .S0 (nx34352)) ;
    aoi22 ix27353 (.Y (nx27352), .A0 (camera_module_cache_ram_75__2), .A1 (
          nx35980), .B0 (camera_module_cache_ram_91__2), .B1 (nx36020)) ;
    dffr camera_module_cache_reg_ram_75__2 (.Q (camera_module_cache_ram_75__2), 
         .QB (\$dummy [721]), .D (nx7153), .CLK (clk), .R (rst)) ;
    mux21_ni ix7154 (.Y (nx7153), .A0 (camera_module_cache_ram_75__2), .A1 (
             nx35266), .S0 (nx34348)) ;
    dffr camera_module_cache_reg_ram_91__2 (.Q (camera_module_cache_ram_91__2), 
         .QB (\$dummy [722]), .D (nx7143), .CLK (clk), .R (rst)) ;
    mux21_ni ix7144 (.Y (nx7143), .A0 (camera_module_cache_ram_91__2), .A1 (
             nx35266), .S0 (nx34344)) ;
    aoi22 ix27361 (.Y (nx27360), .A0 (camera_module_cache_ram_123__2), .A1 (
          nx36060), .B0 (camera_module_cache_ram_107__2), .B1 (nx36100)) ;
    dffr camera_module_cache_reg_ram_123__2 (.Q (camera_module_cache_ram_123__2)
         , .QB (\$dummy [723]), .D (nx7123), .CLK (clk), .R (rst)) ;
    mux21_ni ix7124 (.Y (nx7123), .A0 (camera_module_cache_ram_123__2), .A1 (
             nx35268), .S0 (nx34336)) ;
    dffr camera_module_cache_reg_ram_107__2 (.Q (camera_module_cache_ram_107__2)
         , .QB (\$dummy [724]), .D (nx7133), .CLK (clk), .R (rst)) ;
    mux21_ni ix7134 (.Y (nx7133), .A0 (camera_module_cache_ram_107__2), .A1 (
             nx35268), .S0 (nx34340)) ;
    nand04 ix9607 (.Y (nx9606), .A0 (nx27369), .A1 (nx27377), .A2 (nx27385), .A3 (
           nx27393)) ;
    aoi22 ix27370 (.Y (nx27369), .A0 (camera_module_cache_ram_139__2), .A1 (
          nx36140), .B0 (camera_module_cache_ram_155__2), .B1 (nx36180)) ;
    dffr camera_module_cache_reg_ram_139__2 (.Q (camera_module_cache_ram_139__2)
         , .QB (\$dummy [725]), .D (nx7113), .CLK (clk), .R (rst)) ;
    mux21_ni ix7114 (.Y (nx7113), .A0 (camera_module_cache_ram_139__2), .A1 (
             nx35268), .S0 (nx34332)) ;
    dffr camera_module_cache_reg_ram_155__2 (.Q (camera_module_cache_ram_155__2)
         , .QB (\$dummy [726]), .D (nx7103), .CLK (clk), .R (rst)) ;
    mux21_ni ix7104 (.Y (nx7103), .A0 (camera_module_cache_ram_155__2), .A1 (
             nx35268), .S0 (nx34328)) ;
    aoi22 ix27378 (.Y (nx27377), .A0 (camera_module_cache_ram_187__2), .A1 (
          nx36220), .B0 (camera_module_cache_ram_171__2), .B1 (nx36260)) ;
    dffr camera_module_cache_reg_ram_187__2 (.Q (camera_module_cache_ram_187__2)
         , .QB (\$dummy [727]), .D (nx7083), .CLK (clk), .R (rst)) ;
    mux21_ni ix7084 (.Y (nx7083), .A0 (camera_module_cache_ram_187__2), .A1 (
             nx35268), .S0 (nx34320)) ;
    dffr camera_module_cache_reg_ram_171__2 (.Q (camera_module_cache_ram_171__2)
         , .QB (\$dummy [728]), .D (nx7093), .CLK (clk), .R (rst)) ;
    mux21_ni ix7094 (.Y (nx7093), .A0 (camera_module_cache_ram_171__2), .A1 (
             nx35268), .S0 (nx34324)) ;
    aoi22 ix27386 (.Y (nx27385), .A0 (camera_module_cache_ram_203__2), .A1 (
          nx36300), .B0 (camera_module_cache_ram_219__2), .B1 (nx36340)) ;
    dffr camera_module_cache_reg_ram_203__2 (.Q (camera_module_cache_ram_203__2)
         , .QB (\$dummy [729]), .D (nx7073), .CLK (clk), .R (rst)) ;
    mux21_ni ix7074 (.Y (nx7073), .A0 (camera_module_cache_ram_203__2), .A1 (
             nx35268), .S0 (nx34316)) ;
    dffr camera_module_cache_reg_ram_219__2 (.Q (camera_module_cache_ram_219__2)
         , .QB (\$dummy [730]), .D (nx7063), .CLK (clk), .R (rst)) ;
    mux21_ni ix7064 (.Y (nx7063), .A0 (camera_module_cache_ram_219__2), .A1 (
             nx35270), .S0 (nx34312)) ;
    aoi22 ix27394 (.Y (nx27393), .A0 (camera_module_cache_ram_235__2), .A1 (
          nx36380), .B0 (camera_module_cache_ram_251__2), .B1 (nx36420)) ;
    dffr camera_module_cache_reg_ram_235__2 (.Q (camera_module_cache_ram_235__2)
         , .QB (\$dummy [731]), .D (nx7053), .CLK (clk), .R (rst)) ;
    mux21_ni ix7054 (.Y (nx7053), .A0 (camera_module_cache_ram_235__2), .A1 (
             nx35270), .S0 (nx34308)) ;
    dffr camera_module_cache_reg_ram_251__2 (.Q (camera_module_cache_ram_251__2)
         , .QB (\$dummy [732]), .D (nx7043), .CLK (clk), .R (rst)) ;
    mux21_ni ix7044 (.Y (nx7043), .A0 (camera_module_cache_ram_251__2), .A1 (
             nx35270), .S0 (nx34304)) ;
    nand04 ix9529 (.Y (nx9528), .A0 (nx27402), .A1 (nx27470), .A2 (nx27538), .A3 (
           nx27606)) ;
    oai21 ix27403 (.Y (nx27402), .A0 (nx9518), .A1 (nx9440), .B0 (nx36506)) ;
    nand04 ix9519 (.Y (nx9518), .A0 (nx27405), .A1 (nx27413), .A2 (nx27421), .A3 (
           nx27429)) ;
    aoi22 ix27406 (.Y (nx27405), .A0 (camera_module_cache_ram_12__2), .A1 (
          nx35820), .B0 (camera_module_cache_ram_28__2), .B1 (nx35860)) ;
    dffr camera_module_cache_reg_ram_12__2 (.Q (camera_module_cache_ram_12__2), 
         .QB (\$dummy [733]), .D (nx7033), .CLK (clk), .R (rst)) ;
    mux21_ni ix7034 (.Y (nx7033), .A0 (nx35270), .A1 (
             camera_module_cache_ram_12__2), .S0 (nx36496)) ;
    dffr camera_module_cache_reg_ram_28__2 (.Q (camera_module_cache_ram_28__2), 
         .QB (\$dummy [734]), .D (nx7023), .CLK (clk), .R (rst)) ;
    mux21_ni ix7024 (.Y (nx7023), .A0 (nx35270), .A1 (
             camera_module_cache_ram_28__2), .S0 (nx36510)) ;
    aoi22 ix27414 (.Y (nx27413), .A0 (camera_module_cache_ram_44__2), .A1 (
          nx35900), .B0 (camera_module_cache_ram_60__2), .B1 (nx35940)) ;
    dffr camera_module_cache_reg_ram_44__2 (.Q (camera_module_cache_ram_44__2), 
         .QB (\$dummy [735]), .D (nx7013), .CLK (clk), .R (rst)) ;
    mux21_ni ix7014 (.Y (nx7013), .A0 (nx35270), .A1 (
             camera_module_cache_ram_44__2), .S0 (nx36514)) ;
    dffr camera_module_cache_reg_ram_60__2 (.Q (camera_module_cache_ram_60__2), 
         .QB (\$dummy [736]), .D (nx7003), .CLK (clk), .R (rst)) ;
    mux21_ni ix7004 (.Y (nx7003), .A0 (nx35270), .A1 (
             camera_module_cache_ram_60__2), .S0 (nx36518)) ;
    aoi22 ix27422 (.Y (nx27421), .A0 (camera_module_cache_ram_76__2), .A1 (
          nx35980), .B0 (camera_module_cache_ram_92__2), .B1 (nx36020)) ;
    dffr camera_module_cache_reg_ram_76__2 (.Q (camera_module_cache_ram_76__2), 
         .QB (\$dummy [737]), .D (nx6993), .CLK (clk), .R (rst)) ;
    mux21_ni ix6994 (.Y (nx6993), .A0 (nx35272), .A1 (
             camera_module_cache_ram_76__2), .S0 (nx36522)) ;
    dffr camera_module_cache_reg_ram_92__2 (.Q (camera_module_cache_ram_92__2), 
         .QB (\$dummy [738]), .D (nx6983), .CLK (clk), .R (rst)) ;
    mux21_ni ix6984 (.Y (nx6983), .A0 (nx35272), .A1 (
             camera_module_cache_ram_92__2), .S0 (nx36526)) ;
    aoi22 ix27430 (.Y (nx27429), .A0 (camera_module_cache_ram_124__2), .A1 (
          nx36060), .B0 (camera_module_cache_ram_108__2), .B1 (nx36100)) ;
    dffr camera_module_cache_reg_ram_124__2 (.Q (camera_module_cache_ram_124__2)
         , .QB (\$dummy [739]), .D (nx6963), .CLK (clk), .R (rst)) ;
    mux21_ni ix6964 (.Y (nx6963), .A0 (nx35272), .A1 (
             camera_module_cache_ram_124__2), .S0 (nx36530)) ;
    dffr camera_module_cache_reg_ram_108__2 (.Q (camera_module_cache_ram_108__2)
         , .QB (\$dummy [740]), .D (nx6973), .CLK (clk), .R (rst)) ;
    mux21_ni ix6974 (.Y (nx6973), .A0 (nx35272), .A1 (
             camera_module_cache_ram_108__2), .S0 (nx36534)) ;
    nand04 ix9441 (.Y (nx9440), .A0 (nx27438), .A1 (nx27446), .A2 (nx27454), .A3 (
           nx27462)) ;
    aoi22 ix27439 (.Y (nx27438), .A0 (camera_module_cache_ram_140__2), .A1 (
          nx36140), .B0 (camera_module_cache_ram_156__2), .B1 (nx36180)) ;
    dffr camera_module_cache_reg_ram_140__2 (.Q (camera_module_cache_ram_140__2)
         , .QB (\$dummy [741]), .D (nx6953), .CLK (clk), .R (rst)) ;
    mux21_ni ix6954 (.Y (nx6953), .A0 (nx35272), .A1 (
             camera_module_cache_ram_140__2), .S0 (nx36538)) ;
    dffr camera_module_cache_reg_ram_156__2 (.Q (camera_module_cache_ram_156__2)
         , .QB (\$dummy [742]), .D (nx6943), .CLK (clk), .R (rst)) ;
    mux21_ni ix6944 (.Y (nx6943), .A0 (nx35272), .A1 (
             camera_module_cache_ram_156__2), .S0 (nx36542)) ;
    aoi22 ix27447 (.Y (nx27446), .A0 (camera_module_cache_ram_188__2), .A1 (
          nx36220), .B0 (camera_module_cache_ram_172__2), .B1 (nx36260)) ;
    dffr camera_module_cache_reg_ram_188__2 (.Q (camera_module_cache_ram_188__2)
         , .QB (\$dummy [743]), .D (nx6923), .CLK (clk), .R (rst)) ;
    mux21_ni ix6924 (.Y (nx6923), .A0 (nx35272), .A1 (
             camera_module_cache_ram_188__2), .S0 (nx36546)) ;
    dffr camera_module_cache_reg_ram_172__2 (.Q (camera_module_cache_ram_172__2)
         , .QB (\$dummy [744]), .D (nx6933), .CLK (clk), .R (rst)) ;
    mux21_ni ix6934 (.Y (nx6933), .A0 (nx35274), .A1 (
             camera_module_cache_ram_172__2), .S0 (nx36550)) ;
    aoi22 ix27455 (.Y (nx27454), .A0 (camera_module_cache_ram_204__2), .A1 (
          nx36300), .B0 (camera_module_cache_ram_220__2), .B1 (nx36340)) ;
    dffr camera_module_cache_reg_ram_204__2 (.Q (camera_module_cache_ram_204__2)
         , .QB (\$dummy [745]), .D (nx6913), .CLK (clk), .R (rst)) ;
    mux21_ni ix6914 (.Y (nx6913), .A0 (nx35274), .A1 (
             camera_module_cache_ram_204__2), .S0 (nx36554)) ;
    dffr camera_module_cache_reg_ram_220__2 (.Q (camera_module_cache_ram_220__2)
         , .QB (\$dummy [746]), .D (nx6903), .CLK (clk), .R (rst)) ;
    mux21_ni ix6904 (.Y (nx6903), .A0 (nx35274), .A1 (
             camera_module_cache_ram_220__2), .S0 (nx36558)) ;
    aoi22 ix27463 (.Y (nx27462), .A0 (camera_module_cache_ram_236__2), .A1 (
          nx36380), .B0 (camera_module_cache_ram_252__2), .B1 (nx36420)) ;
    dffr camera_module_cache_reg_ram_236__2 (.Q (camera_module_cache_ram_236__2)
         , .QB (\$dummy [747]), .D (nx6893), .CLK (clk), .R (rst)) ;
    mux21_ni ix6894 (.Y (nx6893), .A0 (nx35274), .A1 (
             camera_module_cache_ram_236__2), .S0 (nx36562)) ;
    dffr camera_module_cache_reg_ram_252__2 (.Q (camera_module_cache_ram_252__2)
         , .QB (\$dummy [748]), .D (nx6883), .CLK (clk), .R (rst)) ;
    mux21_ni ix6884 (.Y (nx6883), .A0 (nx35274), .A1 (
             camera_module_cache_ram_252__2), .S0 (nx36566)) ;
    oai21 ix27471 (.Y (nx27470), .A0 (nx9356), .A1 (nx9278), .B0 (nx36580)) ;
    nand04 ix9357 (.Y (nx9356), .A0 (nx27473), .A1 (nx27481), .A2 (nx27489), .A3 (
           nx27497)) ;
    aoi22 ix27474 (.Y (nx27473), .A0 (camera_module_cache_ram_13__2), .A1 (
          nx35822), .B0 (camera_module_cache_ram_29__2), .B1 (nx35862)) ;
    dffr camera_module_cache_reg_ram_13__2 (.Q (camera_module_cache_ram_13__2), 
         .QB (\$dummy [749]), .D (nx6873), .CLK (clk), .R (rst)) ;
    mux21_ni ix6874 (.Y (nx6873), .A0 (nx35274), .A1 (
             camera_module_cache_ram_13__2), .S0 (nx36570)) ;
    dffr camera_module_cache_reg_ram_29__2 (.Q (camera_module_cache_ram_29__2), 
         .QB (\$dummy [750]), .D (nx6863), .CLK (clk), .R (rst)) ;
    mux21_ni ix6864 (.Y (nx6863), .A0 (nx35274), .A1 (
             camera_module_cache_ram_29__2), .S0 (nx36584)) ;
    aoi22 ix27482 (.Y (nx27481), .A0 (camera_module_cache_ram_45__2), .A1 (
          nx35902), .B0 (camera_module_cache_ram_61__2), .B1 (nx35942)) ;
    dffr camera_module_cache_reg_ram_45__2 (.Q (camera_module_cache_ram_45__2), 
         .QB (\$dummy [751]), .D (nx6853), .CLK (clk), .R (rst)) ;
    mux21_ni ix6854 (.Y (nx6853), .A0 (nx35276), .A1 (
             camera_module_cache_ram_45__2), .S0 (nx36588)) ;
    dffr camera_module_cache_reg_ram_61__2 (.Q (camera_module_cache_ram_61__2), 
         .QB (\$dummy [752]), .D (nx6843), .CLK (clk), .R (rst)) ;
    mux21_ni ix6844 (.Y (nx6843), .A0 (nx35276), .A1 (
             camera_module_cache_ram_61__2), .S0 (nx36592)) ;
    aoi22 ix27490 (.Y (nx27489), .A0 (camera_module_cache_ram_77__2), .A1 (
          nx35982), .B0 (camera_module_cache_ram_93__2), .B1 (nx36022)) ;
    dffr camera_module_cache_reg_ram_77__2 (.Q (camera_module_cache_ram_77__2), 
         .QB (\$dummy [753]), .D (nx6833), .CLK (clk), .R (rst)) ;
    mux21_ni ix6834 (.Y (nx6833), .A0 (nx35276), .A1 (
             camera_module_cache_ram_77__2), .S0 (nx36596)) ;
    dffr camera_module_cache_reg_ram_93__2 (.Q (camera_module_cache_ram_93__2), 
         .QB (\$dummy [754]), .D (nx6823), .CLK (clk), .R (rst)) ;
    mux21_ni ix6824 (.Y (nx6823), .A0 (nx35276), .A1 (
             camera_module_cache_ram_93__2), .S0 (nx36600)) ;
    aoi22 ix27498 (.Y (nx27497), .A0 (camera_module_cache_ram_125__2), .A1 (
          nx36062), .B0 (camera_module_cache_ram_109__2), .B1 (nx36102)) ;
    dffr camera_module_cache_reg_ram_125__2 (.Q (camera_module_cache_ram_125__2)
         , .QB (\$dummy [755]), .D (nx6803), .CLK (clk), .R (rst)) ;
    mux21_ni ix6804 (.Y (nx6803), .A0 (nx35276), .A1 (
             camera_module_cache_ram_125__2), .S0 (nx36604)) ;
    dffr camera_module_cache_reg_ram_109__2 (.Q (camera_module_cache_ram_109__2)
         , .QB (\$dummy [756]), .D (nx6813), .CLK (clk), .R (rst)) ;
    mux21_ni ix6814 (.Y (nx6813), .A0 (nx35276), .A1 (
             camera_module_cache_ram_109__2), .S0 (nx36608)) ;
    nand04 ix9279 (.Y (nx9278), .A0 (nx27506), .A1 (nx27514), .A2 (nx27522), .A3 (
           nx27530)) ;
    aoi22 ix27507 (.Y (nx27506), .A0 (camera_module_cache_ram_141__2), .A1 (
          nx36142), .B0 (camera_module_cache_ram_157__2), .B1 (nx36182)) ;
    dffr camera_module_cache_reg_ram_141__2 (.Q (camera_module_cache_ram_141__2)
         , .QB (\$dummy [757]), .D (nx6793), .CLK (clk), .R (rst)) ;
    mux21_ni ix6794 (.Y (nx6793), .A0 (nx35276), .A1 (
             camera_module_cache_ram_141__2), .S0 (nx36612)) ;
    dffr camera_module_cache_reg_ram_157__2 (.Q (camera_module_cache_ram_157__2)
         , .QB (\$dummy [758]), .D (nx6783), .CLK (clk), .R (rst)) ;
    mux21_ni ix6784 (.Y (nx6783), .A0 (nx35278), .A1 (
             camera_module_cache_ram_157__2), .S0 (nx36616)) ;
    aoi22 ix27515 (.Y (nx27514), .A0 (camera_module_cache_ram_189__2), .A1 (
          nx36222), .B0 (camera_module_cache_ram_173__2), .B1 (nx36262)) ;
    dffr camera_module_cache_reg_ram_189__2 (.Q (camera_module_cache_ram_189__2)
         , .QB (\$dummy [759]), .D (nx6763), .CLK (clk), .R (rst)) ;
    mux21_ni ix6764 (.Y (nx6763), .A0 (nx35278), .A1 (
             camera_module_cache_ram_189__2), .S0 (nx36620)) ;
    dffr camera_module_cache_reg_ram_173__2 (.Q (camera_module_cache_ram_173__2)
         , .QB (\$dummy [760]), .D (nx6773), .CLK (clk), .R (rst)) ;
    mux21_ni ix6774 (.Y (nx6773), .A0 (nx35278), .A1 (
             camera_module_cache_ram_173__2), .S0 (nx36624)) ;
    aoi22 ix27523 (.Y (nx27522), .A0 (camera_module_cache_ram_205__2), .A1 (
          nx36302), .B0 (camera_module_cache_ram_221__2), .B1 (nx36342)) ;
    dffr camera_module_cache_reg_ram_205__2 (.Q (camera_module_cache_ram_205__2)
         , .QB (\$dummy [761]), .D (nx6753), .CLK (clk), .R (rst)) ;
    mux21_ni ix6754 (.Y (nx6753), .A0 (nx35278), .A1 (
             camera_module_cache_ram_205__2), .S0 (nx36628)) ;
    dffr camera_module_cache_reg_ram_221__2 (.Q (camera_module_cache_ram_221__2)
         , .QB (\$dummy [762]), .D (nx6743), .CLK (clk), .R (rst)) ;
    mux21_ni ix6744 (.Y (nx6743), .A0 (nx35278), .A1 (
             camera_module_cache_ram_221__2), .S0 (nx36632)) ;
    aoi22 ix27531 (.Y (nx27530), .A0 (camera_module_cache_ram_237__2), .A1 (
          nx36382), .B0 (camera_module_cache_ram_253__2), .B1 (nx36422)) ;
    dffr camera_module_cache_reg_ram_237__2 (.Q (camera_module_cache_ram_237__2)
         , .QB (\$dummy [763]), .D (nx6733), .CLK (clk), .R (rst)) ;
    mux21_ni ix6734 (.Y (nx6733), .A0 (nx35278), .A1 (
             camera_module_cache_ram_237__2), .S0 (nx36636)) ;
    dffr camera_module_cache_reg_ram_253__2 (.Q (camera_module_cache_ram_253__2)
         , .QB (\$dummy [764]), .D (nx6723), .CLK (clk), .R (rst)) ;
    mux21_ni ix6724 (.Y (nx6723), .A0 (nx35278), .A1 (
             camera_module_cache_ram_253__2), .S0 (nx36640)) ;
    oai21 ix27539 (.Y (nx27538), .A0 (nx9192), .A1 (nx9114), .B0 (nx36654)) ;
    nand04 ix9193 (.Y (nx9192), .A0 (nx27541), .A1 (nx27549), .A2 (nx27557), .A3 (
           nx27565)) ;
    aoi22 ix27542 (.Y (nx27541), .A0 (camera_module_cache_ram_14__2), .A1 (
          nx35822), .B0 (camera_module_cache_ram_30__2), .B1 (nx35862)) ;
    dffr camera_module_cache_reg_ram_14__2 (.Q (camera_module_cache_ram_14__2), 
         .QB (\$dummy [765]), .D (nx6713), .CLK (clk), .R (rst)) ;
    mux21_ni ix6714 (.Y (nx6713), .A0 (nx35280), .A1 (
             camera_module_cache_ram_14__2), .S0 (nx36644)) ;
    dffr camera_module_cache_reg_ram_30__2 (.Q (camera_module_cache_ram_30__2), 
         .QB (\$dummy [766]), .D (nx6703), .CLK (clk), .R (rst)) ;
    mux21_ni ix6704 (.Y (nx6703), .A0 (nx35280), .A1 (
             camera_module_cache_ram_30__2), .S0 (nx36658)) ;
    aoi22 ix27550 (.Y (nx27549), .A0 (camera_module_cache_ram_46__2), .A1 (
          nx35902), .B0 (camera_module_cache_ram_62__2), .B1 (nx35942)) ;
    dffr camera_module_cache_reg_ram_46__2 (.Q (camera_module_cache_ram_46__2), 
         .QB (\$dummy [767]), .D (nx6693), .CLK (clk), .R (rst)) ;
    mux21_ni ix6694 (.Y (nx6693), .A0 (nx35280), .A1 (
             camera_module_cache_ram_46__2), .S0 (nx36662)) ;
    dffr camera_module_cache_reg_ram_62__2 (.Q (camera_module_cache_ram_62__2), 
         .QB (\$dummy [768]), .D (nx6683), .CLK (clk), .R (rst)) ;
    mux21_ni ix6684 (.Y (nx6683), .A0 (nx35280), .A1 (
             camera_module_cache_ram_62__2), .S0 (nx36666)) ;
    aoi22 ix27558 (.Y (nx27557), .A0 (camera_module_cache_ram_78__2), .A1 (
          nx35982), .B0 (camera_module_cache_ram_94__2), .B1 (nx36022)) ;
    dffr camera_module_cache_reg_ram_78__2 (.Q (camera_module_cache_ram_78__2), 
         .QB (\$dummy [769]), .D (nx6673), .CLK (clk), .R (rst)) ;
    mux21_ni ix6674 (.Y (nx6673), .A0 (nx35280), .A1 (
             camera_module_cache_ram_78__2), .S0 (nx36670)) ;
    dffr camera_module_cache_reg_ram_94__2 (.Q (camera_module_cache_ram_94__2), 
         .QB (\$dummy [770]), .D (nx6663), .CLK (clk), .R (rst)) ;
    mux21_ni ix6664 (.Y (nx6663), .A0 (nx35280), .A1 (
             camera_module_cache_ram_94__2), .S0 (nx36674)) ;
    aoi22 ix27566 (.Y (nx27565), .A0 (camera_module_cache_ram_126__2), .A1 (
          nx36062), .B0 (camera_module_cache_ram_110__2), .B1 (nx36102)) ;
    dffr camera_module_cache_reg_ram_126__2 (.Q (camera_module_cache_ram_126__2)
         , .QB (\$dummy [771]), .D (nx6643), .CLK (clk), .R (rst)) ;
    mux21_ni ix6644 (.Y (nx6643), .A0 (nx35280), .A1 (
             camera_module_cache_ram_126__2), .S0 (nx36678)) ;
    dffr camera_module_cache_reg_ram_110__2 (.Q (camera_module_cache_ram_110__2)
         , .QB (\$dummy [772]), .D (nx6653), .CLK (clk), .R (rst)) ;
    mux21_ni ix6654 (.Y (nx6653), .A0 (nx35282), .A1 (
             camera_module_cache_ram_110__2), .S0 (nx36682)) ;
    nand04 ix9115 (.Y (nx9114), .A0 (nx27574), .A1 (nx27582), .A2 (nx27590), .A3 (
           nx27598)) ;
    aoi22 ix27575 (.Y (nx27574), .A0 (camera_module_cache_ram_142__2), .A1 (
          nx36142), .B0 (camera_module_cache_ram_158__2), .B1 (nx36182)) ;
    dffr camera_module_cache_reg_ram_142__2 (.Q (camera_module_cache_ram_142__2)
         , .QB (\$dummy [773]), .D (nx6633), .CLK (clk), .R (rst)) ;
    mux21_ni ix6634 (.Y (nx6633), .A0 (nx35282), .A1 (
             camera_module_cache_ram_142__2), .S0 (nx36686)) ;
    dffr camera_module_cache_reg_ram_158__2 (.Q (camera_module_cache_ram_158__2)
         , .QB (\$dummy [774]), .D (nx6623), .CLK (clk), .R (rst)) ;
    mux21_ni ix6624 (.Y (nx6623), .A0 (nx35282), .A1 (
             camera_module_cache_ram_158__2), .S0 (nx36690)) ;
    aoi22 ix27583 (.Y (nx27582), .A0 (camera_module_cache_ram_190__2), .A1 (
          nx36222), .B0 (camera_module_cache_ram_174__2), .B1 (nx36262)) ;
    dffr camera_module_cache_reg_ram_190__2 (.Q (camera_module_cache_ram_190__2)
         , .QB (\$dummy [775]), .D (nx6603), .CLK (clk), .R (rst)) ;
    mux21_ni ix6604 (.Y (nx6603), .A0 (nx35282), .A1 (
             camera_module_cache_ram_190__2), .S0 (nx36694)) ;
    dffr camera_module_cache_reg_ram_174__2 (.Q (camera_module_cache_ram_174__2)
         , .QB (\$dummy [776]), .D (nx6613), .CLK (clk), .R (rst)) ;
    mux21_ni ix6614 (.Y (nx6613), .A0 (nx35282), .A1 (
             camera_module_cache_ram_174__2), .S0 (nx36698)) ;
    aoi22 ix27591 (.Y (nx27590), .A0 (camera_module_cache_ram_206__2), .A1 (
          nx36302), .B0 (camera_module_cache_ram_222__2), .B1 (nx36342)) ;
    dffr camera_module_cache_reg_ram_206__2 (.Q (camera_module_cache_ram_206__2)
         , .QB (\$dummy [777]), .D (nx6593), .CLK (clk), .R (rst)) ;
    mux21_ni ix6594 (.Y (nx6593), .A0 (nx35282), .A1 (
             camera_module_cache_ram_206__2), .S0 (nx36702)) ;
    dffr camera_module_cache_reg_ram_222__2 (.Q (camera_module_cache_ram_222__2)
         , .QB (\$dummy [778]), .D (nx6583), .CLK (clk), .R (rst)) ;
    mux21_ni ix6584 (.Y (nx6583), .A0 (nx35282), .A1 (
             camera_module_cache_ram_222__2), .S0 (nx36706)) ;
    aoi22 ix27599 (.Y (nx27598), .A0 (camera_module_cache_ram_238__2), .A1 (
          nx36382), .B0 (camera_module_cache_ram_254__2), .B1 (nx36422)) ;
    dffr camera_module_cache_reg_ram_238__2 (.Q (camera_module_cache_ram_238__2)
         , .QB (\$dummy [779]), .D (nx6573), .CLK (clk), .R (rst)) ;
    mux21_ni ix6574 (.Y (nx6573), .A0 (nx35284), .A1 (
             camera_module_cache_ram_238__2), .S0 (nx36710)) ;
    dffr camera_module_cache_reg_ram_254__2 (.Q (camera_module_cache_ram_254__2)
         , .QB (\$dummy [780]), .D (nx6563), .CLK (clk), .R (rst)) ;
    mux21_ni ix6564 (.Y (nx6563), .A0 (nx35284), .A1 (
             camera_module_cache_ram_254__2), .S0 (nx36714)) ;
    oai21 ix27607 (.Y (nx27606), .A0 (nx9030), .A1 (nx8952), .B0 (nx36728)) ;
    nand04 ix9031 (.Y (nx9030), .A0 (nx27609), .A1 (nx27617), .A2 (nx27625), .A3 (
           nx27633)) ;
    aoi22 ix27610 (.Y (nx27609), .A0 (camera_module_cache_ram_15__2), .A1 (
          nx35822), .B0 (camera_module_cache_ram_31__2), .B1 (nx35862)) ;
    dffr camera_module_cache_reg_ram_15__2 (.Q (camera_module_cache_ram_15__2), 
         .QB (\$dummy [781]), .D (nx6553), .CLK (clk), .R (rst)) ;
    mux21_ni ix6554 (.Y (nx6553), .A0 (nx35284), .A1 (
             camera_module_cache_ram_15__2), .S0 (nx36718)) ;
    dffr camera_module_cache_reg_ram_31__2 (.Q (camera_module_cache_ram_31__2), 
         .QB (\$dummy [782]), .D (nx6543), .CLK (clk), .R (rst)) ;
    mux21_ni ix6544 (.Y (nx6543), .A0 (nx35284), .A1 (
             camera_module_cache_ram_31__2), .S0 (nx36732)) ;
    aoi22 ix27618 (.Y (nx27617), .A0 (camera_module_cache_ram_47__2), .A1 (
          nx35902), .B0 (camera_module_cache_ram_63__2), .B1 (nx35942)) ;
    dffr camera_module_cache_reg_ram_47__2 (.Q (camera_module_cache_ram_47__2), 
         .QB (\$dummy [783]), .D (nx6533), .CLK (clk), .R (rst)) ;
    mux21_ni ix6534 (.Y (nx6533), .A0 (nx35284), .A1 (
             camera_module_cache_ram_47__2), .S0 (nx36736)) ;
    dffr camera_module_cache_reg_ram_63__2 (.Q (camera_module_cache_ram_63__2), 
         .QB (\$dummy [784]), .D (nx6523), .CLK (clk), .R (rst)) ;
    mux21_ni ix6524 (.Y (nx6523), .A0 (nx35284), .A1 (
             camera_module_cache_ram_63__2), .S0 (nx36740)) ;
    aoi22 ix27626 (.Y (nx27625), .A0 (camera_module_cache_ram_79__2), .A1 (
          nx35982), .B0 (camera_module_cache_ram_95__2), .B1 (nx36022)) ;
    dffr camera_module_cache_reg_ram_79__2 (.Q (camera_module_cache_ram_79__2), 
         .QB (\$dummy [785]), .D (nx6513), .CLK (clk), .R (rst)) ;
    mux21_ni ix6514 (.Y (nx6513), .A0 (nx35284), .A1 (
             camera_module_cache_ram_79__2), .S0 (nx36744)) ;
    dffr camera_module_cache_reg_ram_95__2 (.Q (camera_module_cache_ram_95__2), 
         .QB (\$dummy [786]), .D (nx6503), .CLK (clk), .R (rst)) ;
    mux21_ni ix6504 (.Y (nx6503), .A0 (nx35286), .A1 (
             camera_module_cache_ram_95__2), .S0 (nx36748)) ;
    aoi22 ix27634 (.Y (nx27633), .A0 (camera_module_cache_ram_127__2), .A1 (
          nx36062), .B0 (camera_module_cache_ram_111__2), .B1 (nx36102)) ;
    dffr camera_module_cache_reg_ram_127__2 (.Q (camera_module_cache_ram_127__2)
         , .QB (\$dummy [787]), .D (nx6483), .CLK (clk), .R (rst)) ;
    mux21_ni ix6484 (.Y (nx6483), .A0 (nx35286), .A1 (
             camera_module_cache_ram_127__2), .S0 (nx36752)) ;
    dffr camera_module_cache_reg_ram_111__2 (.Q (camera_module_cache_ram_111__2)
         , .QB (\$dummy [788]), .D (nx6493), .CLK (clk), .R (rst)) ;
    mux21_ni ix6494 (.Y (nx6493), .A0 (nx35286), .A1 (
             camera_module_cache_ram_111__2), .S0 (nx36756)) ;
    nand04 ix8953 (.Y (nx8952), .A0 (nx27642), .A1 (nx27650), .A2 (nx27658), .A3 (
           nx27666)) ;
    aoi22 ix27643 (.Y (nx27642), .A0 (camera_module_cache_ram_143__2), .A1 (
          nx36142), .B0 (camera_module_cache_ram_159__2), .B1 (nx36182)) ;
    dffr camera_module_cache_reg_ram_143__2 (.Q (camera_module_cache_ram_143__2)
         , .QB (\$dummy [789]), .D (nx6473), .CLK (clk), .R (rst)) ;
    mux21_ni ix6474 (.Y (nx6473), .A0 (nx35286), .A1 (
             camera_module_cache_ram_143__2), .S0 (nx36760)) ;
    dffr camera_module_cache_reg_ram_159__2 (.Q (camera_module_cache_ram_159__2)
         , .QB (\$dummy [790]), .D (nx6463), .CLK (clk), .R (rst)) ;
    mux21_ni ix6464 (.Y (nx6463), .A0 (nx35286), .A1 (
             camera_module_cache_ram_159__2), .S0 (nx36764)) ;
    aoi22 ix27651 (.Y (nx27650), .A0 (camera_module_cache_ram_191__2), .A1 (
          nx36222), .B0 (camera_module_cache_ram_175__2), .B1 (nx36262)) ;
    dffr camera_module_cache_reg_ram_191__2 (.Q (camera_module_cache_ram_191__2)
         , .QB (\$dummy [791]), .D (nx6443), .CLK (clk), .R (rst)) ;
    mux21_ni ix6444 (.Y (nx6443), .A0 (nx35286), .A1 (
             camera_module_cache_ram_191__2), .S0 (nx36768)) ;
    dffr camera_module_cache_reg_ram_175__2 (.Q (camera_module_cache_ram_175__2)
         , .QB (\$dummy [792]), .D (nx6453), .CLK (clk), .R (rst)) ;
    mux21_ni ix6454 (.Y (nx6453), .A0 (nx35286), .A1 (
             camera_module_cache_ram_175__2), .S0 (nx36772)) ;
    aoi22 ix27659 (.Y (nx27658), .A0 (camera_module_cache_ram_207__2), .A1 (
          nx36302), .B0 (camera_module_cache_ram_223__2), .B1 (nx36342)) ;
    dffr camera_module_cache_reg_ram_207__2 (.Q (camera_module_cache_ram_207__2)
         , .QB (\$dummy [793]), .D (nx6433), .CLK (clk), .R (rst)) ;
    mux21_ni ix6434 (.Y (nx6433), .A0 (nx35288), .A1 (
             camera_module_cache_ram_207__2), .S0 (nx36776)) ;
    dffr camera_module_cache_reg_ram_223__2 (.Q (camera_module_cache_ram_223__2)
         , .QB (\$dummy [794]), .D (nx6423), .CLK (clk), .R (rst)) ;
    mux21_ni ix6424 (.Y (nx6423), .A0 (nx35288), .A1 (
             camera_module_cache_ram_223__2), .S0 (nx36780)) ;
    aoi22 ix27667 (.Y (nx27666), .A0 (camera_module_cache_ram_239__2), .A1 (
          nx36382), .B0 (camera_module_cache_ram_255__2), .B1 (nx36422)) ;
    dffr camera_module_cache_reg_ram_239__2 (.Q (camera_module_cache_ram_239__2)
         , .QB (\$dummy [795]), .D (nx6413), .CLK (clk), .R (rst)) ;
    mux21_ni ix6414 (.Y (nx6413), .A0 (nx35288), .A1 (
             camera_module_cache_ram_239__2), .S0 (nx36784)) ;
    dffr camera_module_cache_reg_ram_255__2 (.Q (camera_module_cache_ram_255__2)
         , .QB (\$dummy [796]), .D (nx6403), .CLK (clk), .R (rst)) ;
    mux21_ni ix6404 (.Y (nx6403), .A0 (nx35288), .A1 (
             camera_module_cache_ram_255__2), .S0 (nx36788)) ;
    oai22 ix8755 (.Y (nx8754), .A0 (nx27676), .A1 (nx28817), .B0 (nx29956), .B1 (
          nx8730)) ;
    aoi22 ix27677 (.Y (nx27676), .A0 (camera_module_algo_module_pixel_value_0), 
          .A1 (nx27681), .B0 (one), .B1 (nx5972)) ;
    dff camera_module_algo_module_pixel_reg_reg_q_0 (.Q (
        camera_module_algo_module_pixel_value_0), .QB (\$dummy [797]), .D (
        nx3823), .CLK (clk)) ;
    mux21_ni ix3824 (.Y (nx3823), .A0 (nx5964), .A1 (
             camera_module_algo_module_pixel_value_0), .S0 (nx37152)) ;
    mux21_ni ix27682 (.Y (nx27681), .A0 (nx27683), .A1 (nx35674), .S0 (nx36792)
             ) ;
    nor04 ix27684 (.Y (nx27683), .A0 (nx5944), .A1 (nx4768), .A2 (nx3588), .A3 (
          nx2410)) ;
    nand04 ix5945 (.Y (nx5944), .A0 (nx27686), .A1 (nx27792), .A2 (nx27860), .A3 (
           nx27928)) ;
    oai21 ix27687 (.Y (nx27686), .A0 (nx5934), .A1 (nx5792), .B0 (nx36448)) ;
    nand04 ix5935 (.Y (nx5934), .A0 (nx27689), .A1 (nx27735), .A2 (nx27743), .A3 (
           nx27751)) ;
    aoi22 ix27690 (.Y (nx27689), .A0 (camera_module_cache_ram_0__0), .A1 (
          nx35822), .B0 (camera_module_cache_ram_16__0), .B1 (nx35862)) ;
    dffr camera_module_cache_reg_ram_0__0 (.Q (camera_module_cache_ram_0__0), .QB (
         \$dummy [798]), .D (nx3813), .CLK (clk), .R (rst)) ;
    mux21_ni ix3814 (.Y (nx3813), .A0 (camera_module_cache_ram_0__0), .A1 (
             nx34164), .S0 (nx35134)) ;
    oai221 ix1187 (.Y (nx1186), .A0 (nx34074), .A1 (nx27694), .B0 (nx27710), .B1 (
           nx35712), .C0 (nx27713)) ;
    tri01 nvm_module_tri_dataout_120 (.Y (nvm_data_120), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_112 (.Y (nvm_data_112), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_104 (.Y (nvm_data_104), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_96 (.Y (nvm_data_96), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_88 (.Y (nvm_data_88), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_80 (.Y (nvm_data_80), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_72 (.Y (nvm_data_72), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_64 (.Y (nvm_data_64), .A (nx22549), .E (
          nvm_module_GND0)) ;
    inv01 ix27711 (.Y (nx27710), .A (nvm_data_0)) ;
    tri01 nvm_module_tri_dataout_0 (.Y (nvm_data_0), .A (nx22549), .E (
          nvm_module_GND0)) ;
    nand02 ix27714 (.Y (nx27713), .A0 (nx34074), .A1 (nx1120)) ;
    tri01 nvm_module_tri_dataout_56 (.Y (nvm_data_56), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_48 (.Y (nvm_data_48), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_40 (.Y (nvm_data_40), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_32 (.Y (nvm_data_32), .A (nx22549), .E (
          nvm_module_GND0)) ;
    oai22 ix1089 (.Y (nx1088), .A0 (nx34104), .A1 (nx27724), .B0 (nx34086), .B1 (
          nx27728)) ;
    tri01 nvm_module_tri_dataout_24 (.Y (nvm_data_24), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_16 (.Y (nvm_data_16), .A (nx22549), .E (
          nvm_module_GND0)) ;
    nand02 ix27729 (.Y (nx27728), .A0 (nvm_data_8), .A1 (nx34104)) ;
    tri01 nvm_module_tri_dataout_8 (.Y (nvm_data_8), .A (nx22549), .E (
          nvm_module_GND0)) ;
    dffr camera_module_cache_reg_ram_16__0 (.Q (camera_module_cache_ram_16__0), 
         .QB (\$dummy [799]), .D (nx3803), .CLK (clk), .R (rst)) ;
    mux21_ni ix3804 (.Y (nx3803), .A0 (camera_module_cache_ram_16__0), .A1 (
             nx34164), .S0 (nx35130)) ;
    aoi22 ix27736 (.Y (nx27735), .A0 (camera_module_cache_ram_32__0), .A1 (
          nx35902), .B0 (camera_module_cache_ram_48__0), .B1 (nx35942)) ;
    dffr camera_module_cache_reg_ram_32__0 (.Q (camera_module_cache_ram_32__0), 
         .QB (\$dummy [800]), .D (nx3793), .CLK (clk), .R (rst)) ;
    mux21_ni ix3794 (.Y (nx3793), .A0 (camera_module_cache_ram_32__0), .A1 (
             nx34164), .S0 (nx35126)) ;
    dffr camera_module_cache_reg_ram_48__0 (.Q (camera_module_cache_ram_48__0), 
         .QB (\$dummy [801]), .D (nx3783), .CLK (clk), .R (rst)) ;
    mux21_ni ix3784 (.Y (nx3783), .A0 (camera_module_cache_ram_48__0), .A1 (
             nx34164), .S0 (nx35122)) ;
    aoi22 ix27744 (.Y (nx27743), .A0 (camera_module_cache_ram_64__0), .A1 (
          nx35982), .B0 (camera_module_cache_ram_80__0), .B1 (nx36022)) ;
    dffr camera_module_cache_reg_ram_64__0 (.Q (camera_module_cache_ram_64__0), 
         .QB (\$dummy [802]), .D (nx3773), .CLK (clk), .R (rst)) ;
    mux21_ni ix3774 (.Y (nx3773), .A0 (camera_module_cache_ram_64__0), .A1 (
             nx34164), .S0 (nx35118)) ;
    dffr camera_module_cache_reg_ram_80__0 (.Q (camera_module_cache_ram_80__0), 
         .QB (\$dummy [803]), .D (nx3763), .CLK (clk), .R (rst)) ;
    mux21_ni ix3764 (.Y (nx3763), .A0 (camera_module_cache_ram_80__0), .A1 (
             nx34164), .S0 (nx35114)) ;
    aoi22 ix27752 (.Y (nx27751), .A0 (camera_module_cache_ram_112__0), .A1 (
          nx36062), .B0 (camera_module_cache_ram_96__0), .B1 (nx36102)) ;
    dffr camera_module_cache_reg_ram_112__0 (.Q (camera_module_cache_ram_112__0)
         , .QB (\$dummy [804]), .D (nx3743), .CLK (clk), .R (rst)) ;
    mux21_ni ix3744 (.Y (nx3743), .A0 (camera_module_cache_ram_112__0), .A1 (
             nx34164), .S0 (nx35106)) ;
    dffr camera_module_cache_reg_ram_96__0 (.Q (camera_module_cache_ram_96__0), 
         .QB (\$dummy [805]), .D (nx3753), .CLK (clk), .R (rst)) ;
    mux21_ni ix3754 (.Y (nx3753), .A0 (camera_module_cache_ram_96__0), .A1 (
             nx34166), .S0 (nx35110)) ;
    nand04 ix5793 (.Y (nx5792), .A0 (nx27760), .A1 (nx27768), .A2 (nx27776), .A3 (
           nx27784)) ;
    aoi22 ix27761 (.Y (nx27760), .A0 (camera_module_cache_ram_128__0), .A1 (
          nx36142), .B0 (camera_module_cache_ram_144__0), .B1 (nx36182)) ;
    dffr camera_module_cache_reg_ram_128__0 (.Q (camera_module_cache_ram_128__0)
         , .QB (\$dummy [806]), .D (nx3733), .CLK (clk), .R (rst)) ;
    mux21_ni ix3734 (.Y (nx3733), .A0 (camera_module_cache_ram_128__0), .A1 (
             nx34166), .S0 (nx35102)) ;
    dffr camera_module_cache_reg_ram_144__0 (.Q (camera_module_cache_ram_144__0)
         , .QB (\$dummy [807]), .D (nx3723), .CLK (clk), .R (rst)) ;
    mux21_ni ix3724 (.Y (nx3723), .A0 (camera_module_cache_ram_144__0), .A1 (
             nx34166), .S0 (nx35098)) ;
    aoi22 ix27769 (.Y (nx27768), .A0 (camera_module_cache_ram_176__0), .A1 (
          nx36222), .B0 (camera_module_cache_ram_160__0), .B1 (nx36262)) ;
    dffr camera_module_cache_reg_ram_176__0 (.Q (camera_module_cache_ram_176__0)
         , .QB (\$dummy [808]), .D (nx3703), .CLK (clk), .R (rst)) ;
    mux21_ni ix3704 (.Y (nx3703), .A0 (camera_module_cache_ram_176__0), .A1 (
             nx34166), .S0 (nx35090)) ;
    dffr camera_module_cache_reg_ram_160__0 (.Q (camera_module_cache_ram_160__0)
         , .QB (\$dummy [809]), .D (nx3713), .CLK (clk), .R (rst)) ;
    mux21_ni ix3714 (.Y (nx3713), .A0 (camera_module_cache_ram_160__0), .A1 (
             nx34166), .S0 (nx35094)) ;
    aoi22 ix27777 (.Y (nx27776), .A0 (camera_module_cache_ram_192__0), .A1 (
          nx36302), .B0 (camera_module_cache_ram_208__0), .B1 (nx36342)) ;
    dffr camera_module_cache_reg_ram_192__0 (.Q (camera_module_cache_ram_192__0)
         , .QB (\$dummy [810]), .D (nx3693), .CLK (clk), .R (rst)) ;
    mux21_ni ix3694 (.Y (nx3693), .A0 (camera_module_cache_ram_192__0), .A1 (
             nx34166), .S0 (nx35086)) ;
    dffr camera_module_cache_reg_ram_208__0 (.Q (camera_module_cache_ram_208__0)
         , .QB (\$dummy [811]), .D (nx3683), .CLK (clk), .R (rst)) ;
    mux21_ni ix3684 (.Y (nx3683), .A0 (camera_module_cache_ram_208__0), .A1 (
             nx34166), .S0 (nx35082)) ;
    aoi22 ix27785 (.Y (nx27784), .A0 (camera_module_cache_ram_224__0), .A1 (
          nx36382), .B0 (camera_module_cache_ram_240__0), .B1 (nx36422)) ;
    dffr camera_module_cache_reg_ram_224__0 (.Q (camera_module_cache_ram_224__0)
         , .QB (\$dummy [812]), .D (nx3673), .CLK (clk), .R (rst)) ;
    mux21_ni ix3674 (.Y (nx3673), .A0 (camera_module_cache_ram_224__0), .A1 (
             nx34168), .S0 (nx35078)) ;
    dffr camera_module_cache_reg_ram_240__0 (.Q (camera_module_cache_ram_240__0)
         , .QB (\$dummy [813]), .D (nx3663), .CLK (clk), .R (rst)) ;
    mux21_ni ix3664 (.Y (nx3663), .A0 (camera_module_cache_ram_240__0), .A1 (
             nx34168), .S0 (nx35074)) ;
    oai21 ix27793 (.Y (nx27792), .A0 (nx5642), .A1 (nx5500), .B0 (nx36452)) ;
    nand04 ix5643 (.Y (nx5642), .A0 (nx27795), .A1 (nx27803), .A2 (nx27811), .A3 (
           nx27819)) ;
    aoi22 ix27796 (.Y (nx27795), .A0 (camera_module_cache_ram_1__0), .A1 (
          nx35822), .B0 (camera_module_cache_ram_17__0), .B1 (nx35862)) ;
    dffr camera_module_cache_reg_ram_1__0 (.Q (camera_module_cache_ram_1__0), .QB (
         \$dummy [814]), .D (nx3653), .CLK (clk), .R (rst)) ;
    mux21_ni ix3654 (.Y (nx3653), .A0 (camera_module_cache_ram_1__0), .A1 (
             nx34168), .S0 (nx35064)) ;
    dffr camera_module_cache_reg_ram_17__0 (.Q (camera_module_cache_ram_17__0), 
         .QB (\$dummy [815]), .D (nx3643), .CLK (clk), .R (rst)) ;
    mux21_ni ix3644 (.Y (nx3643), .A0 (camera_module_cache_ram_17__0), .A1 (
             nx34168), .S0 (nx35060)) ;
    aoi22 ix27804 (.Y (nx27803), .A0 (camera_module_cache_ram_33__0), .A1 (
          nx35902), .B0 (camera_module_cache_ram_49__0), .B1 (nx35942)) ;
    dffr camera_module_cache_reg_ram_33__0 (.Q (camera_module_cache_ram_33__0), 
         .QB (\$dummy [816]), .D (nx3633), .CLK (clk), .R (rst)) ;
    mux21_ni ix3634 (.Y (nx3633), .A0 (camera_module_cache_ram_33__0), .A1 (
             nx34168), .S0 (nx35056)) ;
    dffr camera_module_cache_reg_ram_49__0 (.Q (camera_module_cache_ram_49__0), 
         .QB (\$dummy [817]), .D (nx3623), .CLK (clk), .R (rst)) ;
    mux21_ni ix3624 (.Y (nx3623), .A0 (camera_module_cache_ram_49__0), .A1 (
             nx34168), .S0 (nx35052)) ;
    aoi22 ix27812 (.Y (nx27811), .A0 (camera_module_cache_ram_65__0), .A1 (
          nx35982), .B0 (camera_module_cache_ram_81__0), .B1 (nx36022)) ;
    dffr camera_module_cache_reg_ram_65__0 (.Q (camera_module_cache_ram_65__0), 
         .QB (\$dummy [818]), .D (nx3613), .CLK (clk), .R (rst)) ;
    mux21_ni ix3614 (.Y (nx3613), .A0 (camera_module_cache_ram_65__0), .A1 (
             nx34168), .S0 (nx35048)) ;
    dffr camera_module_cache_reg_ram_81__0 (.Q (camera_module_cache_ram_81__0), 
         .QB (\$dummy [819]), .D (nx3603), .CLK (clk), .R (rst)) ;
    mux21_ni ix3604 (.Y (nx3603), .A0 (camera_module_cache_ram_81__0), .A1 (
             nx34170), .S0 (nx35044)) ;
    aoi22 ix27820 (.Y (nx27819), .A0 (camera_module_cache_ram_113__0), .A1 (
          nx36062), .B0 (camera_module_cache_ram_97__0), .B1 (nx36102)) ;
    dffr camera_module_cache_reg_ram_113__0 (.Q (camera_module_cache_ram_113__0)
         , .QB (\$dummy [820]), .D (nx3583), .CLK (clk), .R (rst)) ;
    mux21_ni ix3584 (.Y (nx3583), .A0 (camera_module_cache_ram_113__0), .A1 (
             nx34170), .S0 (nx35036)) ;
    dffr camera_module_cache_reg_ram_97__0 (.Q (camera_module_cache_ram_97__0), 
         .QB (\$dummy [821]), .D (nx3593), .CLK (clk), .R (rst)) ;
    mux21_ni ix3594 (.Y (nx3593), .A0 (camera_module_cache_ram_97__0), .A1 (
             nx34170), .S0 (nx35040)) ;
    nand04 ix5501 (.Y (nx5500), .A0 (nx27828), .A1 (nx27836), .A2 (nx27844), .A3 (
           nx27852)) ;
    aoi22 ix27829 (.Y (nx27828), .A0 (camera_module_cache_ram_129__0), .A1 (
          nx36142), .B0 (camera_module_cache_ram_145__0), .B1 (nx36182)) ;
    dffr camera_module_cache_reg_ram_129__0 (.Q (camera_module_cache_ram_129__0)
         , .QB (\$dummy [822]), .D (nx3573), .CLK (clk), .R (rst)) ;
    mux21_ni ix3574 (.Y (nx3573), .A0 (camera_module_cache_ram_129__0), .A1 (
             nx34170), .S0 (nx35032)) ;
    dffr camera_module_cache_reg_ram_145__0 (.Q (camera_module_cache_ram_145__0)
         , .QB (\$dummy [823]), .D (nx3563), .CLK (clk), .R (rst)) ;
    mux21_ni ix3564 (.Y (nx3563), .A0 (camera_module_cache_ram_145__0), .A1 (
             nx34170), .S0 (nx35028)) ;
    aoi22 ix27837 (.Y (nx27836), .A0 (camera_module_cache_ram_177__0), .A1 (
          nx36222), .B0 (camera_module_cache_ram_161__0), .B1 (nx36262)) ;
    dffr camera_module_cache_reg_ram_177__0 (.Q (camera_module_cache_ram_177__0)
         , .QB (\$dummy [824]), .D (nx3543), .CLK (clk), .R (rst)) ;
    mux21_ni ix3544 (.Y (nx3543), .A0 (camera_module_cache_ram_177__0), .A1 (
             nx34170), .S0 (nx35020)) ;
    dffr camera_module_cache_reg_ram_161__0 (.Q (camera_module_cache_ram_161__0)
         , .QB (\$dummy [825]), .D (nx3553), .CLK (clk), .R (rst)) ;
    mux21_ni ix3554 (.Y (nx3553), .A0 (camera_module_cache_ram_161__0), .A1 (
             nx34170), .S0 (nx35024)) ;
    aoi22 ix27845 (.Y (nx27844), .A0 (camera_module_cache_ram_193__0), .A1 (
          nx36302), .B0 (camera_module_cache_ram_209__0), .B1 (nx36342)) ;
    dffr camera_module_cache_reg_ram_193__0 (.Q (camera_module_cache_ram_193__0)
         , .QB (\$dummy [826]), .D (nx3533), .CLK (clk), .R (rst)) ;
    mux21_ni ix3534 (.Y (nx3533), .A0 (camera_module_cache_ram_193__0), .A1 (
             nx34172), .S0 (nx35016)) ;
    dffr camera_module_cache_reg_ram_209__0 (.Q (camera_module_cache_ram_209__0)
         , .QB (\$dummy [827]), .D (nx3523), .CLK (clk), .R (rst)) ;
    mux21_ni ix3524 (.Y (nx3523), .A0 (camera_module_cache_ram_209__0), .A1 (
             nx34172), .S0 (nx35012)) ;
    aoi22 ix27853 (.Y (nx27852), .A0 (camera_module_cache_ram_225__0), .A1 (
          nx36382), .B0 (camera_module_cache_ram_241__0), .B1 (nx36422)) ;
    dffr camera_module_cache_reg_ram_225__0 (.Q (camera_module_cache_ram_225__0)
         , .QB (\$dummy [828]), .D (nx3513), .CLK (clk), .R (rst)) ;
    mux21_ni ix3514 (.Y (nx3513), .A0 (camera_module_cache_ram_225__0), .A1 (
             nx34172), .S0 (nx35008)) ;
    dffr camera_module_cache_reg_ram_241__0 (.Q (camera_module_cache_ram_241__0)
         , .QB (\$dummy [829]), .D (nx3503), .CLK (clk), .R (rst)) ;
    mux21_ni ix3504 (.Y (nx3503), .A0 (camera_module_cache_ram_241__0), .A1 (
             nx34172), .S0 (nx35004)) ;
    oai21 ix27861 (.Y (nx27860), .A0 (nx5348), .A1 (nx5206), .B0 (nx36456)) ;
    nand04 ix5349 (.Y (nx5348), .A0 (nx27863), .A1 (nx27871), .A2 (nx27879), .A3 (
           nx27887)) ;
    aoi22 ix27864 (.Y (nx27863), .A0 (camera_module_cache_ram_2__0), .A1 (
          nx35822), .B0 (camera_module_cache_ram_18__0), .B1 (nx35862)) ;
    dffr camera_module_cache_reg_ram_2__0 (.Q (camera_module_cache_ram_2__0), .QB (
         \$dummy [830]), .D (nx3493), .CLK (clk), .R (rst)) ;
    mux21_ni ix3494 (.Y (nx3493), .A0 (camera_module_cache_ram_2__0), .A1 (
             nx34172), .S0 (nx34994)) ;
    dffr camera_module_cache_reg_ram_18__0 (.Q (camera_module_cache_ram_18__0), 
         .QB (\$dummy [831]), .D (nx3483), .CLK (clk), .R (rst)) ;
    mux21_ni ix3484 (.Y (nx3483), .A0 (camera_module_cache_ram_18__0), .A1 (
             nx34172), .S0 (nx34990)) ;
    aoi22 ix27872 (.Y (nx27871), .A0 (camera_module_cache_ram_34__0), .A1 (
          nx35902), .B0 (camera_module_cache_ram_50__0), .B1 (nx35942)) ;
    dffr camera_module_cache_reg_ram_34__0 (.Q (camera_module_cache_ram_34__0), 
         .QB (\$dummy [832]), .D (nx3473), .CLK (clk), .R (rst)) ;
    mux21_ni ix3474 (.Y (nx3473), .A0 (camera_module_cache_ram_34__0), .A1 (
             nx34172), .S0 (nx34986)) ;
    dffr camera_module_cache_reg_ram_50__0 (.Q (camera_module_cache_ram_50__0), 
         .QB (\$dummy [833]), .D (nx3463), .CLK (clk), .R (rst)) ;
    mux21_ni ix3464 (.Y (nx3463), .A0 (camera_module_cache_ram_50__0), .A1 (
             nx34174), .S0 (nx34982)) ;
    aoi22 ix27880 (.Y (nx27879), .A0 (camera_module_cache_ram_66__0), .A1 (
          nx35982), .B0 (camera_module_cache_ram_82__0), .B1 (nx36022)) ;
    dffr camera_module_cache_reg_ram_66__0 (.Q (camera_module_cache_ram_66__0), 
         .QB (\$dummy [834]), .D (nx3453), .CLK (clk), .R (rst)) ;
    mux21_ni ix3454 (.Y (nx3453), .A0 (camera_module_cache_ram_66__0), .A1 (
             nx34174), .S0 (nx34978)) ;
    dffr camera_module_cache_reg_ram_82__0 (.Q (camera_module_cache_ram_82__0), 
         .QB (\$dummy [835]), .D (nx3443), .CLK (clk), .R (rst)) ;
    mux21_ni ix3444 (.Y (nx3443), .A0 (camera_module_cache_ram_82__0), .A1 (
             nx34174), .S0 (nx34974)) ;
    aoi22 ix27888 (.Y (nx27887), .A0 (camera_module_cache_ram_114__0), .A1 (
          nx36062), .B0 (camera_module_cache_ram_98__0), .B1 (nx36102)) ;
    dffr camera_module_cache_reg_ram_114__0 (.Q (camera_module_cache_ram_114__0)
         , .QB (\$dummy [836]), .D (nx3423), .CLK (clk), .R (rst)) ;
    mux21_ni ix3424 (.Y (nx3423), .A0 (camera_module_cache_ram_114__0), .A1 (
             nx34174), .S0 (nx34966)) ;
    dffr camera_module_cache_reg_ram_98__0 (.Q (camera_module_cache_ram_98__0), 
         .QB (\$dummy [837]), .D (nx3433), .CLK (clk), .R (rst)) ;
    mux21_ni ix3434 (.Y (nx3433), .A0 (camera_module_cache_ram_98__0), .A1 (
             nx34174), .S0 (nx34970)) ;
    nand04 ix5207 (.Y (nx5206), .A0 (nx27896), .A1 (nx27904), .A2 (nx27912), .A3 (
           nx27920)) ;
    aoi22 ix27897 (.Y (nx27896), .A0 (camera_module_cache_ram_130__0), .A1 (
          nx36142), .B0 (camera_module_cache_ram_146__0), .B1 (nx36182)) ;
    dffr camera_module_cache_reg_ram_130__0 (.Q (camera_module_cache_ram_130__0)
         , .QB (\$dummy [838]), .D (nx3413), .CLK (clk), .R (rst)) ;
    mux21_ni ix3414 (.Y (nx3413), .A0 (camera_module_cache_ram_130__0), .A1 (
             nx34174), .S0 (nx34962)) ;
    dffr camera_module_cache_reg_ram_146__0 (.Q (camera_module_cache_ram_146__0)
         , .QB (\$dummy [839]), .D (nx3403), .CLK (clk), .R (rst)) ;
    mux21_ni ix3404 (.Y (nx3403), .A0 (camera_module_cache_ram_146__0), .A1 (
             nx34174), .S0 (nx34958)) ;
    aoi22 ix27905 (.Y (nx27904), .A0 (camera_module_cache_ram_178__0), .A1 (
          nx36222), .B0 (camera_module_cache_ram_162__0), .B1 (nx36262)) ;
    dffr camera_module_cache_reg_ram_178__0 (.Q (camera_module_cache_ram_178__0)
         , .QB (\$dummy [840]), .D (nx3383), .CLK (clk), .R (rst)) ;
    mux21_ni ix3384 (.Y (nx3383), .A0 (camera_module_cache_ram_178__0), .A1 (
             nx34176), .S0 (nx34950)) ;
    dffr camera_module_cache_reg_ram_162__0 (.Q (camera_module_cache_ram_162__0)
         , .QB (\$dummy [841]), .D (nx3393), .CLK (clk), .R (rst)) ;
    mux21_ni ix3394 (.Y (nx3393), .A0 (camera_module_cache_ram_162__0), .A1 (
             nx34176), .S0 (nx34954)) ;
    aoi22 ix27913 (.Y (nx27912), .A0 (camera_module_cache_ram_194__0), .A1 (
          nx36302), .B0 (camera_module_cache_ram_210__0), .B1 (nx36342)) ;
    dffr camera_module_cache_reg_ram_194__0 (.Q (camera_module_cache_ram_194__0)
         , .QB (\$dummy [842]), .D (nx3373), .CLK (clk), .R (rst)) ;
    mux21_ni ix3374 (.Y (nx3373), .A0 (camera_module_cache_ram_194__0), .A1 (
             nx34176), .S0 (nx34946)) ;
    dffr camera_module_cache_reg_ram_210__0 (.Q (camera_module_cache_ram_210__0)
         , .QB (\$dummy [843]), .D (nx3363), .CLK (clk), .R (rst)) ;
    mux21_ni ix3364 (.Y (nx3363), .A0 (camera_module_cache_ram_210__0), .A1 (
             nx34176), .S0 (nx34942)) ;
    aoi22 ix27921 (.Y (nx27920), .A0 (camera_module_cache_ram_226__0), .A1 (
          nx36382), .B0 (camera_module_cache_ram_242__0), .B1 (nx36422)) ;
    dffr camera_module_cache_reg_ram_226__0 (.Q (camera_module_cache_ram_226__0)
         , .QB (\$dummy [844]), .D (nx3353), .CLK (clk), .R (rst)) ;
    mux21_ni ix3354 (.Y (nx3353), .A0 (camera_module_cache_ram_226__0), .A1 (
             nx34176), .S0 (nx34938)) ;
    dffr camera_module_cache_reg_ram_242__0 (.Q (camera_module_cache_ram_242__0)
         , .QB (\$dummy [845]), .D (nx3343), .CLK (clk), .R (rst)) ;
    mux21_ni ix3344 (.Y (nx3343), .A0 (camera_module_cache_ram_242__0), .A1 (
             nx34176), .S0 (nx34934)) ;
    oai21 ix27929 (.Y (nx27928), .A0 (nx5056), .A1 (nx4914), .B0 (nx36460)) ;
    nand04 ix5057 (.Y (nx5056), .A0 (nx27931), .A1 (nx27939), .A2 (nx27947), .A3 (
           nx27955)) ;
    aoi22 ix27932 (.Y (nx27931), .A0 (camera_module_cache_ram_3__0), .A1 (
          nx35822), .B0 (camera_module_cache_ram_19__0), .B1 (nx35862)) ;
    dffr camera_module_cache_reg_ram_3__0 (.Q (camera_module_cache_ram_3__0), .QB (
         \$dummy [846]), .D (nx3333), .CLK (clk), .R (rst)) ;
    mux21_ni ix3334 (.Y (nx3333), .A0 (camera_module_cache_ram_3__0), .A1 (
             nx34176), .S0 (nx34924)) ;
    dffr camera_module_cache_reg_ram_19__0 (.Q (camera_module_cache_ram_19__0), 
         .QB (\$dummy [847]), .D (nx3323), .CLK (clk), .R (rst)) ;
    mux21_ni ix3324 (.Y (nx3323), .A0 (camera_module_cache_ram_19__0), .A1 (
             nx34178), .S0 (nx34920)) ;
    aoi22 ix27940 (.Y (nx27939), .A0 (camera_module_cache_ram_35__0), .A1 (
          nx35902), .B0 (camera_module_cache_ram_51__0), .B1 (nx35942)) ;
    dffr camera_module_cache_reg_ram_35__0 (.Q (camera_module_cache_ram_35__0), 
         .QB (\$dummy [848]), .D (nx3313), .CLK (clk), .R (rst)) ;
    mux21_ni ix3314 (.Y (nx3313), .A0 (camera_module_cache_ram_35__0), .A1 (
             nx34178), .S0 (nx34916)) ;
    dffr camera_module_cache_reg_ram_51__0 (.Q (camera_module_cache_ram_51__0), 
         .QB (\$dummy [849]), .D (nx3303), .CLK (clk), .R (rst)) ;
    mux21_ni ix3304 (.Y (nx3303), .A0 (camera_module_cache_ram_51__0), .A1 (
             nx34178), .S0 (nx34912)) ;
    aoi22 ix27948 (.Y (nx27947), .A0 (camera_module_cache_ram_67__0), .A1 (
          nx35982), .B0 (camera_module_cache_ram_83__0), .B1 (nx36022)) ;
    dffr camera_module_cache_reg_ram_67__0 (.Q (camera_module_cache_ram_67__0), 
         .QB (\$dummy [850]), .D (nx3293), .CLK (clk), .R (rst)) ;
    mux21_ni ix3294 (.Y (nx3293), .A0 (camera_module_cache_ram_67__0), .A1 (
             nx34178), .S0 (nx34908)) ;
    dffr camera_module_cache_reg_ram_83__0 (.Q (camera_module_cache_ram_83__0), 
         .QB (\$dummy [851]), .D (nx3283), .CLK (clk), .R (rst)) ;
    mux21_ni ix3284 (.Y (nx3283), .A0 (camera_module_cache_ram_83__0), .A1 (
             nx34178), .S0 (nx34904)) ;
    aoi22 ix27956 (.Y (nx27955), .A0 (camera_module_cache_ram_115__0), .A1 (
          nx36062), .B0 (camera_module_cache_ram_99__0), .B1 (nx36102)) ;
    dffr camera_module_cache_reg_ram_115__0 (.Q (camera_module_cache_ram_115__0)
         , .QB (\$dummy [852]), .D (nx3263), .CLK (clk), .R (rst)) ;
    mux21_ni ix3264 (.Y (nx3263), .A0 (camera_module_cache_ram_115__0), .A1 (
             nx34178), .S0 (nx34896)) ;
    dffr camera_module_cache_reg_ram_99__0 (.Q (camera_module_cache_ram_99__0), 
         .QB (\$dummy [853]), .D (nx3273), .CLK (clk), .R (rst)) ;
    mux21_ni ix3274 (.Y (nx3273), .A0 (camera_module_cache_ram_99__0), .A1 (
             nx34178), .S0 (nx34900)) ;
    nand04 ix4915 (.Y (nx4914), .A0 (nx27964), .A1 (nx27972), .A2 (nx27980), .A3 (
           nx27988)) ;
    aoi22 ix27965 (.Y (nx27964), .A0 (camera_module_cache_ram_131__0), .A1 (
          nx36142), .B0 (camera_module_cache_ram_147__0), .B1 (nx36182)) ;
    dffr camera_module_cache_reg_ram_131__0 (.Q (camera_module_cache_ram_131__0)
         , .QB (\$dummy [854]), .D (nx3253), .CLK (clk), .R (rst)) ;
    mux21_ni ix3254 (.Y (nx3253), .A0 (camera_module_cache_ram_131__0), .A1 (
             nx34180), .S0 (nx34892)) ;
    dffr camera_module_cache_reg_ram_147__0 (.Q (camera_module_cache_ram_147__0)
         , .QB (\$dummy [855]), .D (nx3243), .CLK (clk), .R (rst)) ;
    mux21_ni ix3244 (.Y (nx3243), .A0 (camera_module_cache_ram_147__0), .A1 (
             nx34180), .S0 (nx34888)) ;
    aoi22 ix27973 (.Y (nx27972), .A0 (camera_module_cache_ram_179__0), .A1 (
          nx36222), .B0 (camera_module_cache_ram_163__0), .B1 (nx36262)) ;
    dffr camera_module_cache_reg_ram_179__0 (.Q (camera_module_cache_ram_179__0)
         , .QB (\$dummy [856]), .D (nx3223), .CLK (clk), .R (rst)) ;
    mux21_ni ix3224 (.Y (nx3223), .A0 (camera_module_cache_ram_179__0), .A1 (
             nx34180), .S0 (nx34880)) ;
    dffr camera_module_cache_reg_ram_163__0 (.Q (camera_module_cache_ram_163__0)
         , .QB (\$dummy [857]), .D (nx3233), .CLK (clk), .R (rst)) ;
    mux21_ni ix3234 (.Y (nx3233), .A0 (camera_module_cache_ram_163__0), .A1 (
             nx34180), .S0 (nx34884)) ;
    aoi22 ix27981 (.Y (nx27980), .A0 (camera_module_cache_ram_195__0), .A1 (
          nx36302), .B0 (camera_module_cache_ram_211__0), .B1 (nx36342)) ;
    dffr camera_module_cache_reg_ram_195__0 (.Q (camera_module_cache_ram_195__0)
         , .QB (\$dummy [858]), .D (nx3213), .CLK (clk), .R (rst)) ;
    mux21_ni ix3214 (.Y (nx3213), .A0 (camera_module_cache_ram_195__0), .A1 (
             nx34180), .S0 (nx34876)) ;
    dffr camera_module_cache_reg_ram_211__0 (.Q (camera_module_cache_ram_211__0)
         , .QB (\$dummy [859]), .D (nx3203), .CLK (clk), .R (rst)) ;
    mux21_ni ix3204 (.Y (nx3203), .A0 (camera_module_cache_ram_211__0), .A1 (
             nx34180), .S0 (nx34872)) ;
    aoi22 ix27989 (.Y (nx27988), .A0 (camera_module_cache_ram_227__0), .A1 (
          nx36382), .B0 (camera_module_cache_ram_243__0), .B1 (nx36422)) ;
    dffr camera_module_cache_reg_ram_227__0 (.Q (camera_module_cache_ram_227__0)
         , .QB (\$dummy [860]), .D (nx3193), .CLK (clk), .R (rst)) ;
    mux21_ni ix3194 (.Y (nx3193), .A0 (camera_module_cache_ram_227__0), .A1 (
             nx34180), .S0 (nx34868)) ;
    dffr camera_module_cache_reg_ram_243__0 (.Q (camera_module_cache_ram_243__0)
         , .QB (\$dummy [861]), .D (nx3183), .CLK (clk), .R (rst)) ;
    mux21_ni ix3184 (.Y (nx3183), .A0 (camera_module_cache_ram_243__0), .A1 (
             nx34182), .S0 (nx34864)) ;
    nand04 ix4769 (.Y (nx4768), .A0 (nx27997), .A1 (nx28065), .A2 (nx28133), .A3 (
           nx28201)) ;
    oai21 ix27998 (.Y (nx27997), .A0 (nx4758), .A1 (nx4616), .B0 (nx36464)) ;
    nand04 ix4759 (.Y (nx4758), .A0 (nx28000), .A1 (nx28008), .A2 (nx28016), .A3 (
           nx28024)) ;
    aoi22 ix28001 (.Y (nx28000), .A0 (camera_module_cache_ram_4__0), .A1 (
          nx35824), .B0 (camera_module_cache_ram_20__0), .B1 (nx35864)) ;
    dffr camera_module_cache_reg_ram_4__0 (.Q (camera_module_cache_ram_4__0), .QB (
         \$dummy [862]), .D (nx3173), .CLK (clk), .R (rst)) ;
    mux21_ni ix3174 (.Y (nx3173), .A0 (camera_module_cache_ram_4__0), .A1 (
             nx34182), .S0 (nx34854)) ;
    dffr camera_module_cache_reg_ram_20__0 (.Q (camera_module_cache_ram_20__0), 
         .QB (\$dummy [863]), .D (nx3163), .CLK (clk), .R (rst)) ;
    mux21_ni ix3164 (.Y (nx3163), .A0 (camera_module_cache_ram_20__0), .A1 (
             nx34182), .S0 (nx34850)) ;
    aoi22 ix28009 (.Y (nx28008), .A0 (camera_module_cache_ram_36__0), .A1 (
          nx35904), .B0 (camera_module_cache_ram_52__0), .B1 (nx35944)) ;
    dffr camera_module_cache_reg_ram_36__0 (.Q (camera_module_cache_ram_36__0), 
         .QB (\$dummy [864]), .D (nx3153), .CLK (clk), .R (rst)) ;
    mux21_ni ix3154 (.Y (nx3153), .A0 (camera_module_cache_ram_36__0), .A1 (
             nx34182), .S0 (nx34846)) ;
    dffr camera_module_cache_reg_ram_52__0 (.Q (camera_module_cache_ram_52__0), 
         .QB (\$dummy [865]), .D (nx3143), .CLK (clk), .R (rst)) ;
    mux21_ni ix3144 (.Y (nx3143), .A0 (camera_module_cache_ram_52__0), .A1 (
             nx34182), .S0 (nx34842)) ;
    aoi22 ix28017 (.Y (nx28016), .A0 (camera_module_cache_ram_68__0), .A1 (
          nx35984), .B0 (camera_module_cache_ram_84__0), .B1 (nx36024)) ;
    dffr camera_module_cache_reg_ram_68__0 (.Q (camera_module_cache_ram_68__0), 
         .QB (\$dummy [866]), .D (nx3133), .CLK (clk), .R (rst)) ;
    mux21_ni ix3134 (.Y (nx3133), .A0 (camera_module_cache_ram_68__0), .A1 (
             nx34182), .S0 (nx34838)) ;
    dffr camera_module_cache_reg_ram_84__0 (.Q (camera_module_cache_ram_84__0), 
         .QB (\$dummy [867]), .D (nx3123), .CLK (clk), .R (rst)) ;
    mux21_ni ix3124 (.Y (nx3123), .A0 (camera_module_cache_ram_84__0), .A1 (
             nx34182), .S0 (nx34834)) ;
    aoi22 ix28025 (.Y (nx28024), .A0 (camera_module_cache_ram_116__0), .A1 (
          nx36064), .B0 (camera_module_cache_ram_100__0), .B1 (nx36104)) ;
    dffr camera_module_cache_reg_ram_116__0 (.Q (camera_module_cache_ram_116__0)
         , .QB (\$dummy [868]), .D (nx3103), .CLK (clk), .R (rst)) ;
    mux21_ni ix3104 (.Y (nx3103), .A0 (camera_module_cache_ram_116__0), .A1 (
             nx34184), .S0 (nx34826)) ;
    dffr camera_module_cache_reg_ram_100__0 (.Q (camera_module_cache_ram_100__0)
         , .QB (\$dummy [869]), .D (nx3113), .CLK (clk), .R (rst)) ;
    mux21_ni ix3114 (.Y (nx3113), .A0 (camera_module_cache_ram_100__0), .A1 (
             nx34184), .S0 (nx34830)) ;
    nand04 ix4617 (.Y (nx4616), .A0 (nx28033), .A1 (nx28041), .A2 (nx28049), .A3 (
           nx28057)) ;
    aoi22 ix28034 (.Y (nx28033), .A0 (camera_module_cache_ram_132__0), .A1 (
          nx36144), .B0 (camera_module_cache_ram_148__0), .B1 (nx36184)) ;
    dffr camera_module_cache_reg_ram_132__0 (.Q (camera_module_cache_ram_132__0)
         , .QB (\$dummy [870]), .D (nx3093), .CLK (clk), .R (rst)) ;
    mux21_ni ix3094 (.Y (nx3093), .A0 (camera_module_cache_ram_132__0), .A1 (
             nx34184), .S0 (nx34822)) ;
    dffr camera_module_cache_reg_ram_148__0 (.Q (camera_module_cache_ram_148__0)
         , .QB (\$dummy [871]), .D (nx3083), .CLK (clk), .R (rst)) ;
    mux21_ni ix3084 (.Y (nx3083), .A0 (camera_module_cache_ram_148__0), .A1 (
             nx34184), .S0 (nx34818)) ;
    aoi22 ix28042 (.Y (nx28041), .A0 (camera_module_cache_ram_180__0), .A1 (
          nx36224), .B0 (camera_module_cache_ram_164__0), .B1 (nx36264)) ;
    dffr camera_module_cache_reg_ram_180__0 (.Q (camera_module_cache_ram_180__0)
         , .QB (\$dummy [872]), .D (nx3063), .CLK (clk), .R (rst)) ;
    mux21_ni ix3064 (.Y (nx3063), .A0 (camera_module_cache_ram_180__0), .A1 (
             nx34184), .S0 (nx34810)) ;
    dffr camera_module_cache_reg_ram_164__0 (.Q (camera_module_cache_ram_164__0)
         , .QB (\$dummy [873]), .D (nx3073), .CLK (clk), .R (rst)) ;
    mux21_ni ix3074 (.Y (nx3073), .A0 (camera_module_cache_ram_164__0), .A1 (
             nx34184), .S0 (nx34814)) ;
    aoi22 ix28050 (.Y (nx28049), .A0 (camera_module_cache_ram_196__0), .A1 (
          nx36304), .B0 (camera_module_cache_ram_212__0), .B1 (nx36344)) ;
    dffr camera_module_cache_reg_ram_196__0 (.Q (camera_module_cache_ram_196__0)
         , .QB (\$dummy [874]), .D (nx3053), .CLK (clk), .R (rst)) ;
    mux21_ni ix3054 (.Y (nx3053), .A0 (camera_module_cache_ram_196__0), .A1 (
             nx34184), .S0 (nx34806)) ;
    dffr camera_module_cache_reg_ram_212__0 (.Q (camera_module_cache_ram_212__0)
         , .QB (\$dummy [875]), .D (nx3043), .CLK (clk), .R (rst)) ;
    mux21_ni ix3044 (.Y (nx3043), .A0 (camera_module_cache_ram_212__0), .A1 (
             nx34186), .S0 (nx34802)) ;
    aoi22 ix28058 (.Y (nx28057), .A0 (camera_module_cache_ram_228__0), .A1 (
          nx36384), .B0 (camera_module_cache_ram_244__0), .B1 (nx36424)) ;
    dffr camera_module_cache_reg_ram_228__0 (.Q (camera_module_cache_ram_228__0)
         , .QB (\$dummy [876]), .D (nx3033), .CLK (clk), .R (rst)) ;
    mux21_ni ix3034 (.Y (nx3033), .A0 (camera_module_cache_ram_228__0), .A1 (
             nx34186), .S0 (nx34798)) ;
    dffr camera_module_cache_reg_ram_244__0 (.Q (camera_module_cache_ram_244__0)
         , .QB (\$dummy [877]), .D (nx3023), .CLK (clk), .R (rst)) ;
    mux21_ni ix3024 (.Y (nx3023), .A0 (camera_module_cache_ram_244__0), .A1 (
             nx34186), .S0 (nx34794)) ;
    oai21 ix28066 (.Y (nx28065), .A0 (nx4466), .A1 (nx4324), .B0 (nx36468)) ;
    nand04 ix4467 (.Y (nx4466), .A0 (nx28068), .A1 (nx28076), .A2 (nx28084), .A3 (
           nx28092)) ;
    aoi22 ix28069 (.Y (nx28068), .A0 (camera_module_cache_ram_5__0), .A1 (
          nx35824), .B0 (camera_module_cache_ram_21__0), .B1 (nx35864)) ;
    dffr camera_module_cache_reg_ram_5__0 (.Q (camera_module_cache_ram_5__0), .QB (
         \$dummy [878]), .D (nx3013), .CLK (clk), .R (rst)) ;
    mux21_ni ix3014 (.Y (nx3013), .A0 (camera_module_cache_ram_5__0), .A1 (
             nx34186), .S0 (nx34784)) ;
    dffr camera_module_cache_reg_ram_21__0 (.Q (camera_module_cache_ram_21__0), 
         .QB (\$dummy [879]), .D (nx3003), .CLK (clk), .R (rst)) ;
    mux21_ni ix3004 (.Y (nx3003), .A0 (camera_module_cache_ram_21__0), .A1 (
             nx34186), .S0 (nx34780)) ;
    aoi22 ix28077 (.Y (nx28076), .A0 (camera_module_cache_ram_37__0), .A1 (
          nx35904), .B0 (camera_module_cache_ram_53__0), .B1 (nx35944)) ;
    dffr camera_module_cache_reg_ram_37__0 (.Q (camera_module_cache_ram_37__0), 
         .QB (\$dummy [880]), .D (nx2993), .CLK (clk), .R (rst)) ;
    mux21_ni ix2994 (.Y (nx2993), .A0 (camera_module_cache_ram_37__0), .A1 (
             nx34186), .S0 (nx34776)) ;
    dffr camera_module_cache_reg_ram_53__0 (.Q (camera_module_cache_ram_53__0), 
         .QB (\$dummy [881]), .D (nx2983), .CLK (clk), .R (rst)) ;
    mux21_ni ix2984 (.Y (nx2983), .A0 (camera_module_cache_ram_53__0), .A1 (
             nx34186), .S0 (nx34772)) ;
    aoi22 ix28085 (.Y (nx28084), .A0 (camera_module_cache_ram_69__0), .A1 (
          nx35984), .B0 (camera_module_cache_ram_85__0), .B1 (nx36024)) ;
    dffr camera_module_cache_reg_ram_69__0 (.Q (camera_module_cache_ram_69__0), 
         .QB (\$dummy [882]), .D (nx2973), .CLK (clk), .R (rst)) ;
    mux21_ni ix2974 (.Y (nx2973), .A0 (camera_module_cache_ram_69__0), .A1 (
             nx34188), .S0 (nx34768)) ;
    dffr camera_module_cache_reg_ram_85__0 (.Q (camera_module_cache_ram_85__0), 
         .QB (\$dummy [883]), .D (nx2963), .CLK (clk), .R (rst)) ;
    mux21_ni ix2964 (.Y (nx2963), .A0 (camera_module_cache_ram_85__0), .A1 (
             nx34188), .S0 (nx34764)) ;
    aoi22 ix28093 (.Y (nx28092), .A0 (camera_module_cache_ram_117__0), .A1 (
          nx36064), .B0 (camera_module_cache_ram_101__0), .B1 (nx36104)) ;
    dffr camera_module_cache_reg_ram_117__0 (.Q (camera_module_cache_ram_117__0)
         , .QB (\$dummy [884]), .D (nx2943), .CLK (clk), .R (rst)) ;
    mux21_ni ix2944 (.Y (nx2943), .A0 (camera_module_cache_ram_117__0), .A1 (
             nx34188), .S0 (nx34756)) ;
    dffr camera_module_cache_reg_ram_101__0 (.Q (camera_module_cache_ram_101__0)
         , .QB (\$dummy [885]), .D (nx2953), .CLK (clk), .R (rst)) ;
    mux21_ni ix2954 (.Y (nx2953), .A0 (camera_module_cache_ram_101__0), .A1 (
             nx34188), .S0 (nx34760)) ;
    nand04 ix4325 (.Y (nx4324), .A0 (nx28101), .A1 (nx28109), .A2 (nx28117), .A3 (
           nx28125)) ;
    aoi22 ix28102 (.Y (nx28101), .A0 (camera_module_cache_ram_133__0), .A1 (
          nx36144), .B0 (camera_module_cache_ram_149__0), .B1 (nx36184)) ;
    dffr camera_module_cache_reg_ram_133__0 (.Q (camera_module_cache_ram_133__0)
         , .QB (\$dummy [886]), .D (nx2933), .CLK (clk), .R (rst)) ;
    mux21_ni ix2934 (.Y (nx2933), .A0 (camera_module_cache_ram_133__0), .A1 (
             nx34188), .S0 (nx34752)) ;
    dffr camera_module_cache_reg_ram_149__0 (.Q (camera_module_cache_ram_149__0)
         , .QB (\$dummy [887]), .D (nx2923), .CLK (clk), .R (rst)) ;
    mux21_ni ix2924 (.Y (nx2923), .A0 (camera_module_cache_ram_149__0), .A1 (
             nx34188), .S0 (nx34748)) ;
    aoi22 ix28110 (.Y (nx28109), .A0 (camera_module_cache_ram_181__0), .A1 (
          nx36224), .B0 (camera_module_cache_ram_165__0), .B1 (nx36264)) ;
    dffr camera_module_cache_reg_ram_181__0 (.Q (camera_module_cache_ram_181__0)
         , .QB (\$dummy [888]), .D (nx2903), .CLK (clk), .R (rst)) ;
    mux21_ni ix2904 (.Y (nx2903), .A0 (camera_module_cache_ram_181__0), .A1 (
             nx34188), .S0 (nx34740)) ;
    dffr camera_module_cache_reg_ram_165__0 (.Q (camera_module_cache_ram_165__0)
         , .QB (\$dummy [889]), .D (nx2913), .CLK (clk), .R (rst)) ;
    mux21_ni ix2914 (.Y (nx2913), .A0 (camera_module_cache_ram_165__0), .A1 (
             nx34190), .S0 (nx34744)) ;
    aoi22 ix28118 (.Y (nx28117), .A0 (camera_module_cache_ram_197__0), .A1 (
          nx36304), .B0 (camera_module_cache_ram_213__0), .B1 (nx36344)) ;
    dffr camera_module_cache_reg_ram_197__0 (.Q (camera_module_cache_ram_197__0)
         , .QB (\$dummy [890]), .D (nx2893), .CLK (clk), .R (rst)) ;
    mux21_ni ix2894 (.Y (nx2893), .A0 (camera_module_cache_ram_197__0), .A1 (
             nx34190), .S0 (nx34736)) ;
    dffr camera_module_cache_reg_ram_213__0 (.Q (camera_module_cache_ram_213__0)
         , .QB (\$dummy [891]), .D (nx2883), .CLK (clk), .R (rst)) ;
    mux21_ni ix2884 (.Y (nx2883), .A0 (camera_module_cache_ram_213__0), .A1 (
             nx34190), .S0 (nx34732)) ;
    aoi22 ix28126 (.Y (nx28125), .A0 (camera_module_cache_ram_229__0), .A1 (
          nx36384), .B0 (camera_module_cache_ram_245__0), .B1 (nx36424)) ;
    dffr camera_module_cache_reg_ram_229__0 (.Q (camera_module_cache_ram_229__0)
         , .QB (\$dummy [892]), .D (nx2873), .CLK (clk), .R (rst)) ;
    mux21_ni ix2874 (.Y (nx2873), .A0 (camera_module_cache_ram_229__0), .A1 (
             nx34190), .S0 (nx34728)) ;
    dffr camera_module_cache_reg_ram_245__0 (.Q (camera_module_cache_ram_245__0)
         , .QB (\$dummy [893]), .D (nx2863), .CLK (clk), .R (rst)) ;
    mux21_ni ix2864 (.Y (nx2863), .A0 (camera_module_cache_ram_245__0), .A1 (
             nx34190), .S0 (nx34724)) ;
    oai21 ix28134 (.Y (nx28133), .A0 (nx4172), .A1 (nx4030), .B0 (nx36472)) ;
    nand04 ix4173 (.Y (nx4172), .A0 (nx28136), .A1 (nx28144), .A2 (nx28152), .A3 (
           nx28160)) ;
    aoi22 ix28137 (.Y (nx28136), .A0 (camera_module_cache_ram_6__0), .A1 (
          nx35824), .B0 (camera_module_cache_ram_22__0), .B1 (nx35864)) ;
    dffr camera_module_cache_reg_ram_6__0 (.Q (camera_module_cache_ram_6__0), .QB (
         \$dummy [894]), .D (nx2853), .CLK (clk), .R (rst)) ;
    mux21_ni ix2854 (.Y (nx2853), .A0 (camera_module_cache_ram_6__0), .A1 (
             nx34190), .S0 (nx34714)) ;
    dffr camera_module_cache_reg_ram_22__0 (.Q (camera_module_cache_ram_22__0), 
         .QB (\$dummy [895]), .D (nx2843), .CLK (clk), .R (rst)) ;
    mux21_ni ix2844 (.Y (nx2843), .A0 (camera_module_cache_ram_22__0), .A1 (
             nx34190), .S0 (nx34710)) ;
    aoi22 ix28145 (.Y (nx28144), .A0 (camera_module_cache_ram_38__0), .A1 (
          nx35904), .B0 (camera_module_cache_ram_54__0), .B1 (nx35944)) ;
    dffr camera_module_cache_reg_ram_38__0 (.Q (camera_module_cache_ram_38__0), 
         .QB (\$dummy [896]), .D (nx2833), .CLK (clk), .R (rst)) ;
    mux21_ni ix2834 (.Y (nx2833), .A0 (camera_module_cache_ram_38__0), .A1 (
             nx34192), .S0 (nx34706)) ;
    dffr camera_module_cache_reg_ram_54__0 (.Q (camera_module_cache_ram_54__0), 
         .QB (\$dummy [897]), .D (nx2823), .CLK (clk), .R (rst)) ;
    mux21_ni ix2824 (.Y (nx2823), .A0 (camera_module_cache_ram_54__0), .A1 (
             nx34192), .S0 (nx34702)) ;
    aoi22 ix28153 (.Y (nx28152), .A0 (camera_module_cache_ram_70__0), .A1 (
          nx35984), .B0 (camera_module_cache_ram_86__0), .B1 (nx36024)) ;
    dffr camera_module_cache_reg_ram_70__0 (.Q (camera_module_cache_ram_70__0), 
         .QB (\$dummy [898]), .D (nx2813), .CLK (clk), .R (rst)) ;
    mux21_ni ix2814 (.Y (nx2813), .A0 (camera_module_cache_ram_70__0), .A1 (
             nx34192), .S0 (nx34698)) ;
    dffr camera_module_cache_reg_ram_86__0 (.Q (camera_module_cache_ram_86__0), 
         .QB (\$dummy [899]), .D (nx2803), .CLK (clk), .R (rst)) ;
    mux21_ni ix2804 (.Y (nx2803), .A0 (camera_module_cache_ram_86__0), .A1 (
             nx34192), .S0 (nx34694)) ;
    aoi22 ix28161 (.Y (nx28160), .A0 (camera_module_cache_ram_118__0), .A1 (
          nx36064), .B0 (camera_module_cache_ram_102__0), .B1 (nx36104)) ;
    dffr camera_module_cache_reg_ram_118__0 (.Q (camera_module_cache_ram_118__0)
         , .QB (\$dummy [900]), .D (nx2783), .CLK (clk), .R (rst)) ;
    mux21_ni ix2784 (.Y (nx2783), .A0 (camera_module_cache_ram_118__0), .A1 (
             nx34192), .S0 (nx34686)) ;
    dffr camera_module_cache_reg_ram_102__0 (.Q (camera_module_cache_ram_102__0)
         , .QB (\$dummy [901]), .D (nx2793), .CLK (clk), .R (rst)) ;
    mux21_ni ix2794 (.Y (nx2793), .A0 (camera_module_cache_ram_102__0), .A1 (
             nx34192), .S0 (nx34690)) ;
    nand04 ix4031 (.Y (nx4030), .A0 (nx28169), .A1 (nx28177), .A2 (nx28185), .A3 (
           nx28193)) ;
    aoi22 ix28170 (.Y (nx28169), .A0 (camera_module_cache_ram_134__0), .A1 (
          nx36144), .B0 (camera_module_cache_ram_150__0), .B1 (nx36184)) ;
    dffr camera_module_cache_reg_ram_134__0 (.Q (camera_module_cache_ram_134__0)
         , .QB (\$dummy [902]), .D (nx2773), .CLK (clk), .R (rst)) ;
    mux21_ni ix2774 (.Y (nx2773), .A0 (camera_module_cache_ram_134__0), .A1 (
             nx34192), .S0 (nx34682)) ;
    dffr camera_module_cache_reg_ram_150__0 (.Q (camera_module_cache_ram_150__0)
         , .QB (\$dummy [903]), .D (nx2763), .CLK (clk), .R (rst)) ;
    mux21_ni ix2764 (.Y (nx2763), .A0 (camera_module_cache_ram_150__0), .A1 (
             nx34194), .S0 (nx34678)) ;
    aoi22 ix28178 (.Y (nx28177), .A0 (camera_module_cache_ram_182__0), .A1 (
          nx36224), .B0 (camera_module_cache_ram_166__0), .B1 (nx36264)) ;
    dffr camera_module_cache_reg_ram_182__0 (.Q (camera_module_cache_ram_182__0)
         , .QB (\$dummy [904]), .D (nx2743), .CLK (clk), .R (rst)) ;
    mux21_ni ix2744 (.Y (nx2743), .A0 (camera_module_cache_ram_182__0), .A1 (
             nx34194), .S0 (nx34670)) ;
    dffr camera_module_cache_reg_ram_166__0 (.Q (camera_module_cache_ram_166__0)
         , .QB (\$dummy [905]), .D (nx2753), .CLK (clk), .R (rst)) ;
    mux21_ni ix2754 (.Y (nx2753), .A0 (camera_module_cache_ram_166__0), .A1 (
             nx34194), .S0 (nx34674)) ;
    aoi22 ix28186 (.Y (nx28185), .A0 (camera_module_cache_ram_198__0), .A1 (
          nx36304), .B0 (camera_module_cache_ram_214__0), .B1 (nx36344)) ;
    dffr camera_module_cache_reg_ram_198__0 (.Q (camera_module_cache_ram_198__0)
         , .QB (\$dummy [906]), .D (nx2733), .CLK (clk), .R (rst)) ;
    mux21_ni ix2734 (.Y (nx2733), .A0 (camera_module_cache_ram_198__0), .A1 (
             nx34194), .S0 (nx34666)) ;
    dffr camera_module_cache_reg_ram_214__0 (.Q (camera_module_cache_ram_214__0)
         , .QB (\$dummy [907]), .D (nx2723), .CLK (clk), .R (rst)) ;
    mux21_ni ix2724 (.Y (nx2723), .A0 (camera_module_cache_ram_214__0), .A1 (
             nx34194), .S0 (nx34662)) ;
    aoi22 ix28194 (.Y (nx28193), .A0 (camera_module_cache_ram_230__0), .A1 (
          nx36384), .B0 (camera_module_cache_ram_246__0), .B1 (nx36424)) ;
    dffr camera_module_cache_reg_ram_230__0 (.Q (camera_module_cache_ram_230__0)
         , .QB (\$dummy [908]), .D (nx2713), .CLK (clk), .R (rst)) ;
    mux21_ni ix2714 (.Y (nx2713), .A0 (camera_module_cache_ram_230__0), .A1 (
             nx34194), .S0 (nx34658)) ;
    dffr camera_module_cache_reg_ram_246__0 (.Q (camera_module_cache_ram_246__0)
         , .QB (\$dummy [909]), .D (nx2703), .CLK (clk), .R (rst)) ;
    mux21_ni ix2704 (.Y (nx2703), .A0 (camera_module_cache_ram_246__0), .A1 (
             nx34194), .S0 (nx34654)) ;
    oai21 ix28202 (.Y (nx28201), .A0 (nx3880), .A1 (nx3738), .B0 (nx36476)) ;
    nand04 ix3881 (.Y (nx3880), .A0 (nx28204), .A1 (nx28212), .A2 (nx28220), .A3 (
           nx28228)) ;
    aoi22 ix28205 (.Y (nx28204), .A0 (camera_module_cache_ram_7__0), .A1 (
          nx35824), .B0 (camera_module_cache_ram_23__0), .B1 (nx35864)) ;
    dffr camera_module_cache_reg_ram_7__0 (.Q (camera_module_cache_ram_7__0), .QB (
         \$dummy [910]), .D (nx2693), .CLK (clk), .R (rst)) ;
    mux21_ni ix2694 (.Y (nx2693), .A0 (camera_module_cache_ram_7__0), .A1 (
             nx34196), .S0 (nx34644)) ;
    dffr camera_module_cache_reg_ram_23__0 (.Q (camera_module_cache_ram_23__0), 
         .QB (\$dummy [911]), .D (nx2683), .CLK (clk), .R (rst)) ;
    mux21_ni ix2684 (.Y (nx2683), .A0 (camera_module_cache_ram_23__0), .A1 (
             nx34196), .S0 (nx34640)) ;
    aoi22 ix28213 (.Y (nx28212), .A0 (camera_module_cache_ram_39__0), .A1 (
          nx35904), .B0 (camera_module_cache_ram_55__0), .B1 (nx35944)) ;
    dffr camera_module_cache_reg_ram_39__0 (.Q (camera_module_cache_ram_39__0), 
         .QB (\$dummy [912]), .D (nx2673), .CLK (clk), .R (rst)) ;
    mux21_ni ix2674 (.Y (nx2673), .A0 (camera_module_cache_ram_39__0), .A1 (
             nx34196), .S0 (nx34636)) ;
    dffr camera_module_cache_reg_ram_55__0 (.Q (camera_module_cache_ram_55__0), 
         .QB (\$dummy [913]), .D (nx2663), .CLK (clk), .R (rst)) ;
    mux21_ni ix2664 (.Y (nx2663), .A0 (camera_module_cache_ram_55__0), .A1 (
             nx34196), .S0 (nx34632)) ;
    aoi22 ix28221 (.Y (nx28220), .A0 (camera_module_cache_ram_71__0), .A1 (
          nx35984), .B0 (camera_module_cache_ram_87__0), .B1 (nx36024)) ;
    dffr camera_module_cache_reg_ram_71__0 (.Q (camera_module_cache_ram_71__0), 
         .QB (\$dummy [914]), .D (nx2653), .CLK (clk), .R (rst)) ;
    mux21_ni ix2654 (.Y (nx2653), .A0 (camera_module_cache_ram_71__0), .A1 (
             nx34196), .S0 (nx34628)) ;
    dffr camera_module_cache_reg_ram_87__0 (.Q (camera_module_cache_ram_87__0), 
         .QB (\$dummy [915]), .D (nx2643), .CLK (clk), .R (rst)) ;
    mux21_ni ix2644 (.Y (nx2643), .A0 (camera_module_cache_ram_87__0), .A1 (
             nx34196), .S0 (nx34624)) ;
    aoi22 ix28229 (.Y (nx28228), .A0 (camera_module_cache_ram_119__0), .A1 (
          nx36064), .B0 (camera_module_cache_ram_103__0), .B1 (nx36104)) ;
    dffr camera_module_cache_reg_ram_119__0 (.Q (camera_module_cache_ram_119__0)
         , .QB (\$dummy [916]), .D (nx2623), .CLK (clk), .R (rst)) ;
    mux21_ni ix2624 (.Y (nx2623), .A0 (camera_module_cache_ram_119__0), .A1 (
             nx34196), .S0 (nx34616)) ;
    dffr camera_module_cache_reg_ram_103__0 (.Q (camera_module_cache_ram_103__0)
         , .QB (\$dummy [917]), .D (nx2633), .CLK (clk), .R (rst)) ;
    mux21_ni ix2634 (.Y (nx2633), .A0 (camera_module_cache_ram_103__0), .A1 (
             nx34198), .S0 (nx34620)) ;
    nand04 ix3739 (.Y (nx3738), .A0 (nx28237), .A1 (nx28245), .A2 (nx28253), .A3 (
           nx28261)) ;
    aoi22 ix28238 (.Y (nx28237), .A0 (camera_module_cache_ram_135__0), .A1 (
          nx36144), .B0 (camera_module_cache_ram_151__0), .B1 (nx36184)) ;
    dffr camera_module_cache_reg_ram_135__0 (.Q (camera_module_cache_ram_135__0)
         , .QB (\$dummy [918]), .D (nx2613), .CLK (clk), .R (rst)) ;
    mux21_ni ix2614 (.Y (nx2613), .A0 (camera_module_cache_ram_135__0), .A1 (
             nx34198), .S0 (nx34612)) ;
    dffr camera_module_cache_reg_ram_151__0 (.Q (camera_module_cache_ram_151__0)
         , .QB (\$dummy [919]), .D (nx2603), .CLK (clk), .R (rst)) ;
    mux21_ni ix2604 (.Y (nx2603), .A0 (camera_module_cache_ram_151__0), .A1 (
             nx34198), .S0 (nx34608)) ;
    aoi22 ix28246 (.Y (nx28245), .A0 (camera_module_cache_ram_183__0), .A1 (
          nx36224), .B0 (camera_module_cache_ram_167__0), .B1 (nx36264)) ;
    dffr camera_module_cache_reg_ram_183__0 (.Q (camera_module_cache_ram_183__0)
         , .QB (\$dummy [920]), .D (nx2583), .CLK (clk), .R (rst)) ;
    mux21_ni ix2584 (.Y (nx2583), .A0 (camera_module_cache_ram_183__0), .A1 (
             nx34198), .S0 (nx34600)) ;
    dffr camera_module_cache_reg_ram_167__0 (.Q (camera_module_cache_ram_167__0)
         , .QB (\$dummy [921]), .D (nx2593), .CLK (clk), .R (rst)) ;
    mux21_ni ix2594 (.Y (nx2593), .A0 (camera_module_cache_ram_167__0), .A1 (
             nx34198), .S0 (nx34604)) ;
    aoi22 ix28254 (.Y (nx28253), .A0 (camera_module_cache_ram_199__0), .A1 (
          nx36304), .B0 (camera_module_cache_ram_215__0), .B1 (nx36344)) ;
    dffr camera_module_cache_reg_ram_199__0 (.Q (camera_module_cache_ram_199__0)
         , .QB (\$dummy [922]), .D (nx2573), .CLK (clk), .R (rst)) ;
    mux21_ni ix2574 (.Y (nx2573), .A0 (camera_module_cache_ram_199__0), .A1 (
             nx34198), .S0 (nx34596)) ;
    dffr camera_module_cache_reg_ram_215__0 (.Q (camera_module_cache_ram_215__0)
         , .QB (\$dummy [923]), .D (nx2563), .CLK (clk), .R (rst)) ;
    mux21_ni ix2564 (.Y (nx2563), .A0 (camera_module_cache_ram_215__0), .A1 (
             nx34198), .S0 (nx34592)) ;
    aoi22 ix28262 (.Y (nx28261), .A0 (camera_module_cache_ram_231__0), .A1 (
          nx36384), .B0 (camera_module_cache_ram_247__0), .B1 (nx36424)) ;
    dffr camera_module_cache_reg_ram_231__0 (.Q (camera_module_cache_ram_231__0)
         , .QB (\$dummy [924]), .D (nx2553), .CLK (clk), .R (rst)) ;
    mux21_ni ix2554 (.Y (nx2553), .A0 (camera_module_cache_ram_231__0), .A1 (
             nx34200), .S0 (nx34588)) ;
    dffr camera_module_cache_reg_ram_247__0 (.Q (camera_module_cache_ram_247__0)
         , .QB (\$dummy [925]), .D (nx2543), .CLK (clk), .R (rst)) ;
    mux21_ni ix2544 (.Y (nx2543), .A0 (camera_module_cache_ram_247__0), .A1 (
             nx34200), .S0 (nx34584)) ;
    nand04 ix3589 (.Y (nx3588), .A0 (nx28270), .A1 (nx28338), .A2 (nx28406), .A3 (
           nx28474)) ;
    oai21 ix28271 (.Y (nx28270), .A0 (nx3578), .A1 (nx3436), .B0 (nx36480)) ;
    nand04 ix3579 (.Y (nx3578), .A0 (nx28273), .A1 (nx28281), .A2 (nx28289), .A3 (
           nx28297)) ;
    aoi22 ix28274 (.Y (nx28273), .A0 (camera_module_cache_ram_8__0), .A1 (
          nx35824), .B0 (camera_module_cache_ram_24__0), .B1 (nx35864)) ;
    dffr camera_module_cache_reg_ram_8__0 (.Q (camera_module_cache_ram_8__0), .QB (
         \$dummy [926]), .D (nx2533), .CLK (clk), .R (rst)) ;
    mux21_ni ix2534 (.Y (nx2533), .A0 (camera_module_cache_ram_8__0), .A1 (
             nx34200), .S0 (nx34574)) ;
    dffr camera_module_cache_reg_ram_24__0 (.Q (camera_module_cache_ram_24__0), 
         .QB (\$dummy [927]), .D (nx2523), .CLK (clk), .R (rst)) ;
    mux21_ni ix2524 (.Y (nx2523), .A0 (camera_module_cache_ram_24__0), .A1 (
             nx34200), .S0 (nx34570)) ;
    aoi22 ix28282 (.Y (nx28281), .A0 (camera_module_cache_ram_40__0), .A1 (
          nx35904), .B0 (camera_module_cache_ram_56__0), .B1 (nx35944)) ;
    dffr camera_module_cache_reg_ram_40__0 (.Q (camera_module_cache_ram_40__0), 
         .QB (\$dummy [928]), .D (nx2513), .CLK (clk), .R (rst)) ;
    mux21_ni ix2514 (.Y (nx2513), .A0 (camera_module_cache_ram_40__0), .A1 (
             nx34200), .S0 (nx34566)) ;
    dffr camera_module_cache_reg_ram_56__0 (.Q (camera_module_cache_ram_56__0), 
         .QB (\$dummy [929]), .D (nx2503), .CLK (clk), .R (rst)) ;
    mux21_ni ix2504 (.Y (nx2503), .A0 (camera_module_cache_ram_56__0), .A1 (
             nx34200), .S0 (nx34562)) ;
    aoi22 ix28290 (.Y (nx28289), .A0 (camera_module_cache_ram_72__0), .A1 (
          nx35984), .B0 (camera_module_cache_ram_88__0), .B1 (nx36024)) ;
    dffr camera_module_cache_reg_ram_72__0 (.Q (camera_module_cache_ram_72__0), 
         .QB (\$dummy [930]), .D (nx2493), .CLK (clk), .R (rst)) ;
    mux21_ni ix2494 (.Y (nx2493), .A0 (camera_module_cache_ram_72__0), .A1 (
             nx34200), .S0 (nx34558)) ;
    dffr camera_module_cache_reg_ram_88__0 (.Q (camera_module_cache_ram_88__0), 
         .QB (\$dummy [931]), .D (nx2483), .CLK (clk), .R (rst)) ;
    mux21_ni ix2484 (.Y (nx2483), .A0 (camera_module_cache_ram_88__0), .A1 (
             nx34202), .S0 (nx34554)) ;
    aoi22 ix28298 (.Y (nx28297), .A0 (camera_module_cache_ram_120__0), .A1 (
          nx36064), .B0 (camera_module_cache_ram_104__0), .B1 (nx36104)) ;
    dffr camera_module_cache_reg_ram_120__0 (.Q (camera_module_cache_ram_120__0)
         , .QB (\$dummy [932]), .D (nx2463), .CLK (clk), .R (rst)) ;
    mux21_ni ix2464 (.Y (nx2463), .A0 (camera_module_cache_ram_120__0), .A1 (
             nx34202), .S0 (nx34546)) ;
    dffr camera_module_cache_reg_ram_104__0 (.Q (camera_module_cache_ram_104__0)
         , .QB (\$dummy [933]), .D (nx2473), .CLK (clk), .R (rst)) ;
    mux21_ni ix2474 (.Y (nx2473), .A0 (camera_module_cache_ram_104__0), .A1 (
             nx34202), .S0 (nx34550)) ;
    nand04 ix3437 (.Y (nx3436), .A0 (nx28306), .A1 (nx28314), .A2 (nx28322), .A3 (
           nx28330)) ;
    aoi22 ix28307 (.Y (nx28306), .A0 (camera_module_cache_ram_136__0), .A1 (
          nx36144), .B0 (camera_module_cache_ram_152__0), .B1 (nx36184)) ;
    dffr camera_module_cache_reg_ram_136__0 (.Q (camera_module_cache_ram_136__0)
         , .QB (\$dummy [934]), .D (nx2453), .CLK (clk), .R (rst)) ;
    mux21_ni ix2454 (.Y (nx2453), .A0 (camera_module_cache_ram_136__0), .A1 (
             nx34202), .S0 (nx34542)) ;
    dffr camera_module_cache_reg_ram_152__0 (.Q (camera_module_cache_ram_152__0)
         , .QB (\$dummy [935]), .D (nx2443), .CLK (clk), .R (rst)) ;
    mux21_ni ix2444 (.Y (nx2443), .A0 (camera_module_cache_ram_152__0), .A1 (
             nx34202), .S0 (nx34538)) ;
    aoi22 ix28315 (.Y (nx28314), .A0 (camera_module_cache_ram_184__0), .A1 (
          nx36224), .B0 (camera_module_cache_ram_168__0), .B1 (nx36264)) ;
    dffr camera_module_cache_reg_ram_184__0 (.Q (camera_module_cache_ram_184__0)
         , .QB (\$dummy [936]), .D (nx2423), .CLK (clk), .R (rst)) ;
    mux21_ni ix2424 (.Y (nx2423), .A0 (camera_module_cache_ram_184__0), .A1 (
             nx34202), .S0 (nx34530)) ;
    dffr camera_module_cache_reg_ram_168__0 (.Q (camera_module_cache_ram_168__0)
         , .QB (\$dummy [937]), .D (nx2433), .CLK (clk), .R (rst)) ;
    mux21_ni ix2434 (.Y (nx2433), .A0 (camera_module_cache_ram_168__0), .A1 (
             nx34202), .S0 (nx34534)) ;
    aoi22 ix28323 (.Y (nx28322), .A0 (camera_module_cache_ram_200__0), .A1 (
          nx36304), .B0 (camera_module_cache_ram_216__0), .B1 (nx36344)) ;
    dffr camera_module_cache_reg_ram_200__0 (.Q (camera_module_cache_ram_200__0)
         , .QB (\$dummy [938]), .D (nx2413), .CLK (clk), .R (rst)) ;
    mux21_ni ix2414 (.Y (nx2413), .A0 (camera_module_cache_ram_200__0), .A1 (
             nx34204), .S0 (nx34526)) ;
    dffr camera_module_cache_reg_ram_216__0 (.Q (camera_module_cache_ram_216__0)
         , .QB (\$dummy [939]), .D (nx2403), .CLK (clk), .R (rst)) ;
    mux21_ni ix2404 (.Y (nx2403), .A0 (camera_module_cache_ram_216__0), .A1 (
             nx34204), .S0 (nx34522)) ;
    aoi22 ix28331 (.Y (nx28330), .A0 (camera_module_cache_ram_232__0), .A1 (
          nx36384), .B0 (camera_module_cache_ram_248__0), .B1 (nx36424)) ;
    dffr camera_module_cache_reg_ram_232__0 (.Q (camera_module_cache_ram_232__0)
         , .QB (\$dummy [940]), .D (nx2393), .CLK (clk), .R (rst)) ;
    mux21_ni ix2394 (.Y (nx2393), .A0 (camera_module_cache_ram_232__0), .A1 (
             nx34204), .S0 (nx34518)) ;
    dffr camera_module_cache_reg_ram_248__0 (.Q (camera_module_cache_ram_248__0)
         , .QB (\$dummy [941]), .D (nx2383), .CLK (clk), .R (rst)) ;
    mux21_ni ix2384 (.Y (nx2383), .A0 (camera_module_cache_ram_248__0), .A1 (
             nx34204), .S0 (nx34514)) ;
    oai21 ix28339 (.Y (nx28338), .A0 (nx3286), .A1 (nx3144), .B0 (nx36484)) ;
    nand04 ix3287 (.Y (nx3286), .A0 (nx28341), .A1 (nx28349), .A2 (nx28357), .A3 (
           nx28365)) ;
    aoi22 ix28342 (.Y (nx28341), .A0 (camera_module_cache_ram_9__0), .A1 (
          nx35824), .B0 (camera_module_cache_ram_25__0), .B1 (nx35864)) ;
    dffr camera_module_cache_reg_ram_9__0 (.Q (camera_module_cache_ram_9__0), .QB (
         \$dummy [942]), .D (nx2373), .CLK (clk), .R (rst)) ;
    mux21_ni ix2374 (.Y (nx2373), .A0 (camera_module_cache_ram_9__0), .A1 (
             nx34204), .S0 (nx34504)) ;
    dffr camera_module_cache_reg_ram_25__0 (.Q (camera_module_cache_ram_25__0), 
         .QB (\$dummy [943]), .D (nx2363), .CLK (clk), .R (rst)) ;
    mux21_ni ix2364 (.Y (nx2363), .A0 (camera_module_cache_ram_25__0), .A1 (
             nx34204), .S0 (nx34500)) ;
    aoi22 ix28350 (.Y (nx28349), .A0 (camera_module_cache_ram_41__0), .A1 (
          nx35904), .B0 (camera_module_cache_ram_57__0), .B1 (nx35944)) ;
    dffr camera_module_cache_reg_ram_41__0 (.Q (camera_module_cache_ram_41__0), 
         .QB (\$dummy [944]), .D (nx2353), .CLK (clk), .R (rst)) ;
    mux21_ni ix2354 (.Y (nx2353), .A0 (camera_module_cache_ram_41__0), .A1 (
             nx34204), .S0 (nx34496)) ;
    dffr camera_module_cache_reg_ram_57__0 (.Q (camera_module_cache_ram_57__0), 
         .QB (\$dummy [945]), .D (nx2343), .CLK (clk), .R (rst)) ;
    mux21_ni ix2344 (.Y (nx2343), .A0 (camera_module_cache_ram_57__0), .A1 (
             nx34206), .S0 (nx34492)) ;
    aoi22 ix28358 (.Y (nx28357), .A0 (camera_module_cache_ram_73__0), .A1 (
          nx35984), .B0 (camera_module_cache_ram_89__0), .B1 (nx36024)) ;
    dffr camera_module_cache_reg_ram_73__0 (.Q (camera_module_cache_ram_73__0), 
         .QB (\$dummy [946]), .D (nx2333), .CLK (clk), .R (rst)) ;
    mux21_ni ix2334 (.Y (nx2333), .A0 (camera_module_cache_ram_73__0), .A1 (
             nx34206), .S0 (nx34488)) ;
    dffr camera_module_cache_reg_ram_89__0 (.Q (camera_module_cache_ram_89__0), 
         .QB (\$dummy [947]), .D (nx2323), .CLK (clk), .R (rst)) ;
    mux21_ni ix2324 (.Y (nx2323), .A0 (camera_module_cache_ram_89__0), .A1 (
             nx34206), .S0 (nx34484)) ;
    aoi22 ix28366 (.Y (nx28365), .A0 (camera_module_cache_ram_121__0), .A1 (
          nx36064), .B0 (camera_module_cache_ram_105__0), .B1 (nx36104)) ;
    dffr camera_module_cache_reg_ram_121__0 (.Q (camera_module_cache_ram_121__0)
         , .QB (\$dummy [948]), .D (nx2303), .CLK (clk), .R (rst)) ;
    mux21_ni ix2304 (.Y (nx2303), .A0 (camera_module_cache_ram_121__0), .A1 (
             nx34206), .S0 (nx34476)) ;
    dffr camera_module_cache_reg_ram_105__0 (.Q (camera_module_cache_ram_105__0)
         , .QB (\$dummy [949]), .D (nx2313), .CLK (clk), .R (rst)) ;
    mux21_ni ix2314 (.Y (nx2313), .A0 (camera_module_cache_ram_105__0), .A1 (
             nx34206), .S0 (nx34480)) ;
    nand04 ix3145 (.Y (nx3144), .A0 (nx28374), .A1 (nx28382), .A2 (nx28390), .A3 (
           nx28398)) ;
    aoi22 ix28375 (.Y (nx28374), .A0 (camera_module_cache_ram_137__0), .A1 (
          nx36144), .B0 (camera_module_cache_ram_153__0), .B1 (nx36184)) ;
    dffr camera_module_cache_reg_ram_137__0 (.Q (camera_module_cache_ram_137__0)
         , .QB (\$dummy [950]), .D (nx2293), .CLK (clk), .R (rst)) ;
    mux21_ni ix2294 (.Y (nx2293), .A0 (camera_module_cache_ram_137__0), .A1 (
             nx34206), .S0 (nx34472)) ;
    dffr camera_module_cache_reg_ram_153__0 (.Q (camera_module_cache_ram_153__0)
         , .QB (\$dummy [951]), .D (nx2283), .CLK (clk), .R (rst)) ;
    mux21_ni ix2284 (.Y (nx2283), .A0 (camera_module_cache_ram_153__0), .A1 (
             nx34206), .S0 (nx34468)) ;
    aoi22 ix28383 (.Y (nx28382), .A0 (camera_module_cache_ram_185__0), .A1 (
          nx36224), .B0 (camera_module_cache_ram_169__0), .B1 (nx36264)) ;
    dffr camera_module_cache_reg_ram_185__0 (.Q (camera_module_cache_ram_185__0)
         , .QB (\$dummy [952]), .D (nx2263), .CLK (clk), .R (rst)) ;
    mux21_ni ix2264 (.Y (nx2263), .A0 (camera_module_cache_ram_185__0), .A1 (
             nx34208), .S0 (nx34460)) ;
    dffr camera_module_cache_reg_ram_169__0 (.Q (camera_module_cache_ram_169__0)
         , .QB (\$dummy [953]), .D (nx2273), .CLK (clk), .R (rst)) ;
    mux21_ni ix2274 (.Y (nx2273), .A0 (camera_module_cache_ram_169__0), .A1 (
             nx34208), .S0 (nx34464)) ;
    aoi22 ix28391 (.Y (nx28390), .A0 (camera_module_cache_ram_201__0), .A1 (
          nx36304), .B0 (camera_module_cache_ram_217__0), .B1 (nx36344)) ;
    dffr camera_module_cache_reg_ram_201__0 (.Q (camera_module_cache_ram_201__0)
         , .QB (\$dummy [954]), .D (nx2253), .CLK (clk), .R (rst)) ;
    mux21_ni ix2254 (.Y (nx2253), .A0 (camera_module_cache_ram_201__0), .A1 (
             nx34208), .S0 (nx34456)) ;
    dffr camera_module_cache_reg_ram_217__0 (.Q (camera_module_cache_ram_217__0)
         , .QB (\$dummy [955]), .D (nx2243), .CLK (clk), .R (rst)) ;
    mux21_ni ix2244 (.Y (nx2243), .A0 (camera_module_cache_ram_217__0), .A1 (
             nx34208), .S0 (nx34452)) ;
    aoi22 ix28399 (.Y (nx28398), .A0 (camera_module_cache_ram_233__0), .A1 (
          nx36384), .B0 (camera_module_cache_ram_249__0), .B1 (nx36424)) ;
    dffr camera_module_cache_reg_ram_233__0 (.Q (camera_module_cache_ram_233__0)
         , .QB (\$dummy [956]), .D (nx2233), .CLK (clk), .R (rst)) ;
    mux21_ni ix2234 (.Y (nx2233), .A0 (camera_module_cache_ram_233__0), .A1 (
             nx34208), .S0 (nx34448)) ;
    dffr camera_module_cache_reg_ram_249__0 (.Q (camera_module_cache_ram_249__0)
         , .QB (\$dummy [957]), .D (nx2223), .CLK (clk), .R (rst)) ;
    mux21_ni ix2224 (.Y (nx2223), .A0 (camera_module_cache_ram_249__0), .A1 (
             nx34208), .S0 (nx34444)) ;
    oai21 ix28407 (.Y (nx28406), .A0 (nx2992), .A1 (nx2850), .B0 (nx36488)) ;
    nand04 ix2993 (.Y (nx2992), .A0 (nx28409), .A1 (nx28417), .A2 (nx28425), .A3 (
           nx28433)) ;
    aoi22 ix28410 (.Y (nx28409), .A0 (camera_module_cache_ram_10__0), .A1 (
          nx35824), .B0 (camera_module_cache_ram_26__0), .B1 (nx35864)) ;
    dffr camera_module_cache_reg_ram_10__0 (.Q (camera_module_cache_ram_10__0), 
         .QB (\$dummy [958]), .D (nx2213), .CLK (clk), .R (rst)) ;
    mux21_ni ix2214 (.Y (nx2213), .A0 (camera_module_cache_ram_10__0), .A1 (
             nx34208), .S0 (nx34434)) ;
    dffr camera_module_cache_reg_ram_26__0 (.Q (camera_module_cache_ram_26__0), 
         .QB (\$dummy [959]), .D (nx2203), .CLK (clk), .R (rst)) ;
    mux21_ni ix2204 (.Y (nx2203), .A0 (camera_module_cache_ram_26__0), .A1 (
             nx34210), .S0 (nx34430)) ;
    aoi22 ix28418 (.Y (nx28417), .A0 (camera_module_cache_ram_42__0), .A1 (
          nx35904), .B0 (camera_module_cache_ram_58__0), .B1 (nx35944)) ;
    dffr camera_module_cache_reg_ram_42__0 (.Q (camera_module_cache_ram_42__0), 
         .QB (\$dummy [960]), .D (nx2193), .CLK (clk), .R (rst)) ;
    mux21_ni ix2194 (.Y (nx2193), .A0 (camera_module_cache_ram_42__0), .A1 (
             nx34210), .S0 (nx34426)) ;
    dffr camera_module_cache_reg_ram_58__0 (.Q (camera_module_cache_ram_58__0), 
         .QB (\$dummy [961]), .D (nx2183), .CLK (clk), .R (rst)) ;
    mux21_ni ix2184 (.Y (nx2183), .A0 (camera_module_cache_ram_58__0), .A1 (
             nx34210), .S0 (nx34422)) ;
    aoi22 ix28426 (.Y (nx28425), .A0 (camera_module_cache_ram_74__0), .A1 (
          nx35984), .B0 (camera_module_cache_ram_90__0), .B1 (nx36024)) ;
    dffr camera_module_cache_reg_ram_74__0 (.Q (camera_module_cache_ram_74__0), 
         .QB (\$dummy [962]), .D (nx2173), .CLK (clk), .R (rst)) ;
    mux21_ni ix2174 (.Y (nx2173), .A0 (camera_module_cache_ram_74__0), .A1 (
             nx34210), .S0 (nx34418)) ;
    dffr camera_module_cache_reg_ram_90__0 (.Q (camera_module_cache_ram_90__0), 
         .QB (\$dummy [963]), .D (nx2163), .CLK (clk), .R (rst)) ;
    mux21_ni ix2164 (.Y (nx2163), .A0 (camera_module_cache_ram_90__0), .A1 (
             nx34210), .S0 (nx34414)) ;
    aoi22 ix28434 (.Y (nx28433), .A0 (camera_module_cache_ram_122__0), .A1 (
          nx36064), .B0 (camera_module_cache_ram_106__0), .B1 (nx36104)) ;
    dffr camera_module_cache_reg_ram_122__0 (.Q (camera_module_cache_ram_122__0)
         , .QB (\$dummy [964]), .D (nx2143), .CLK (clk), .R (rst)) ;
    mux21_ni ix2144 (.Y (nx2143), .A0 (camera_module_cache_ram_122__0), .A1 (
             nx34210), .S0 (nx34406)) ;
    dffr camera_module_cache_reg_ram_106__0 (.Q (camera_module_cache_ram_106__0)
         , .QB (\$dummy [965]), .D (nx2153), .CLK (clk), .R (rst)) ;
    mux21_ni ix2154 (.Y (nx2153), .A0 (camera_module_cache_ram_106__0), .A1 (
             nx34210), .S0 (nx34410)) ;
    nand04 ix2851 (.Y (nx2850), .A0 (nx28442), .A1 (nx28450), .A2 (nx28458), .A3 (
           nx28466)) ;
    aoi22 ix28443 (.Y (nx28442), .A0 (camera_module_cache_ram_138__0), .A1 (
          nx36144), .B0 (camera_module_cache_ram_154__0), .B1 (nx36184)) ;
    dffr camera_module_cache_reg_ram_138__0 (.Q (camera_module_cache_ram_138__0)
         , .QB (\$dummy [966]), .D (nx2133), .CLK (clk), .R (rst)) ;
    mux21_ni ix2134 (.Y (nx2133), .A0 (camera_module_cache_ram_138__0), .A1 (
             nx34212), .S0 (nx34402)) ;
    dffr camera_module_cache_reg_ram_154__0 (.Q (camera_module_cache_ram_154__0)
         , .QB (\$dummy [967]), .D (nx2123), .CLK (clk), .R (rst)) ;
    mux21_ni ix2124 (.Y (nx2123), .A0 (camera_module_cache_ram_154__0), .A1 (
             nx34212), .S0 (nx34398)) ;
    aoi22 ix28451 (.Y (nx28450), .A0 (camera_module_cache_ram_186__0), .A1 (
          nx36224), .B0 (camera_module_cache_ram_170__0), .B1 (nx36264)) ;
    dffr camera_module_cache_reg_ram_186__0 (.Q (camera_module_cache_ram_186__0)
         , .QB (\$dummy [968]), .D (nx2103), .CLK (clk), .R (rst)) ;
    mux21_ni ix2104 (.Y (nx2103), .A0 (camera_module_cache_ram_186__0), .A1 (
             nx34212), .S0 (nx34390)) ;
    dffr camera_module_cache_reg_ram_170__0 (.Q (camera_module_cache_ram_170__0)
         , .QB (\$dummy [969]), .D (nx2113), .CLK (clk), .R (rst)) ;
    mux21_ni ix2114 (.Y (nx2113), .A0 (camera_module_cache_ram_170__0), .A1 (
             nx34212), .S0 (nx34394)) ;
    aoi22 ix28459 (.Y (nx28458), .A0 (camera_module_cache_ram_202__0), .A1 (
          nx36304), .B0 (camera_module_cache_ram_218__0), .B1 (nx36344)) ;
    dffr camera_module_cache_reg_ram_202__0 (.Q (camera_module_cache_ram_202__0)
         , .QB (\$dummy [970]), .D (nx2093), .CLK (clk), .R (rst)) ;
    mux21_ni ix2094 (.Y (nx2093), .A0 (camera_module_cache_ram_202__0), .A1 (
             nx34212), .S0 (nx34386)) ;
    dffr camera_module_cache_reg_ram_218__0 (.Q (camera_module_cache_ram_218__0)
         , .QB (\$dummy [971]), .D (nx2083), .CLK (clk), .R (rst)) ;
    mux21_ni ix2084 (.Y (nx2083), .A0 (camera_module_cache_ram_218__0), .A1 (
             nx34212), .S0 (nx34382)) ;
    aoi22 ix28467 (.Y (nx28466), .A0 (camera_module_cache_ram_234__0), .A1 (
          nx36384), .B0 (camera_module_cache_ram_250__0), .B1 (nx36424)) ;
    dffr camera_module_cache_reg_ram_234__0 (.Q (camera_module_cache_ram_234__0)
         , .QB (\$dummy [972]), .D (nx2073), .CLK (clk), .R (rst)) ;
    mux21_ni ix2074 (.Y (nx2073), .A0 (camera_module_cache_ram_234__0), .A1 (
             nx34212), .S0 (nx34378)) ;
    dffr camera_module_cache_reg_ram_250__0 (.Q (camera_module_cache_ram_250__0)
         , .QB (\$dummy [973]), .D (nx2063), .CLK (clk), .R (rst)) ;
    mux21_ni ix2064 (.Y (nx2063), .A0 (camera_module_cache_ram_250__0), .A1 (
             nx34214), .S0 (nx34374)) ;
    oai21 ix28475 (.Y (nx28474), .A0 (nx2700), .A1 (nx2558), .B0 (nx36492)) ;
    nand04 ix2701 (.Y (nx2700), .A0 (nx28477), .A1 (nx28485), .A2 (nx28493), .A3 (
           nx28501)) ;
    aoi22 ix28478 (.Y (nx28477), .A0 (camera_module_cache_ram_11__0), .A1 (
          nx35826), .B0 (camera_module_cache_ram_27__0), .B1 (nx35866)) ;
    dffr camera_module_cache_reg_ram_11__0 (.Q (camera_module_cache_ram_11__0), 
         .QB (\$dummy [974]), .D (nx2053), .CLK (clk), .R (rst)) ;
    mux21_ni ix2054 (.Y (nx2053), .A0 (camera_module_cache_ram_11__0), .A1 (
             nx34214), .S0 (nx34364)) ;
    dffr camera_module_cache_reg_ram_27__0 (.Q (camera_module_cache_ram_27__0), 
         .QB (\$dummy [975]), .D (nx2043), .CLK (clk), .R (rst)) ;
    mux21_ni ix2044 (.Y (nx2043), .A0 (camera_module_cache_ram_27__0), .A1 (
             nx34214), .S0 (nx34360)) ;
    aoi22 ix28486 (.Y (nx28485), .A0 (camera_module_cache_ram_43__0), .A1 (
          nx35906), .B0 (camera_module_cache_ram_59__0), .B1 (nx35946)) ;
    dffr camera_module_cache_reg_ram_43__0 (.Q (camera_module_cache_ram_43__0), 
         .QB (\$dummy [976]), .D (nx2033), .CLK (clk), .R (rst)) ;
    mux21_ni ix2034 (.Y (nx2033), .A0 (camera_module_cache_ram_43__0), .A1 (
             nx34214), .S0 (nx34356)) ;
    dffr camera_module_cache_reg_ram_59__0 (.Q (camera_module_cache_ram_59__0), 
         .QB (\$dummy [977]), .D (nx2023), .CLK (clk), .R (rst)) ;
    mux21_ni ix2024 (.Y (nx2023), .A0 (camera_module_cache_ram_59__0), .A1 (
             nx34214), .S0 (nx34352)) ;
    aoi22 ix28494 (.Y (nx28493), .A0 (camera_module_cache_ram_75__0), .A1 (
          nx35986), .B0 (camera_module_cache_ram_91__0), .B1 (nx36026)) ;
    dffr camera_module_cache_reg_ram_75__0 (.Q (camera_module_cache_ram_75__0), 
         .QB (\$dummy [978]), .D (nx2013), .CLK (clk), .R (rst)) ;
    mux21_ni ix2014 (.Y (nx2013), .A0 (camera_module_cache_ram_75__0), .A1 (
             nx34214), .S0 (nx34348)) ;
    dffr camera_module_cache_reg_ram_91__0 (.Q (camera_module_cache_ram_91__0), 
         .QB (\$dummy [979]), .D (nx2003), .CLK (clk), .R (rst)) ;
    mux21_ni ix2004 (.Y (nx2003), .A0 (camera_module_cache_ram_91__0), .A1 (
             nx34214), .S0 (nx34344)) ;
    aoi22 ix28502 (.Y (nx28501), .A0 (camera_module_cache_ram_123__0), .A1 (
          nx36066), .B0 (camera_module_cache_ram_107__0), .B1 (nx36106)) ;
    dffr camera_module_cache_reg_ram_123__0 (.Q (camera_module_cache_ram_123__0)
         , .QB (\$dummy [980]), .D (nx1983), .CLK (clk), .R (rst)) ;
    mux21_ni ix1984 (.Y (nx1983), .A0 (camera_module_cache_ram_123__0), .A1 (
             nx34216), .S0 (nx34336)) ;
    dffr camera_module_cache_reg_ram_107__0 (.Q (camera_module_cache_ram_107__0)
         , .QB (\$dummy [981]), .D (nx1993), .CLK (clk), .R (rst)) ;
    mux21_ni ix1994 (.Y (nx1993), .A0 (camera_module_cache_ram_107__0), .A1 (
             nx34216), .S0 (nx34340)) ;
    nand04 ix2559 (.Y (nx2558), .A0 (nx28510), .A1 (nx28518), .A2 (nx28526), .A3 (
           nx28534)) ;
    aoi22 ix28511 (.Y (nx28510), .A0 (camera_module_cache_ram_139__0), .A1 (
          nx36146), .B0 (camera_module_cache_ram_155__0), .B1 (nx36186)) ;
    dffr camera_module_cache_reg_ram_139__0 (.Q (camera_module_cache_ram_139__0)
         , .QB (\$dummy [982]), .D (nx1973), .CLK (clk), .R (rst)) ;
    mux21_ni ix1974 (.Y (nx1973), .A0 (camera_module_cache_ram_139__0), .A1 (
             nx34216), .S0 (nx34332)) ;
    dffr camera_module_cache_reg_ram_155__0 (.Q (camera_module_cache_ram_155__0)
         , .QB (\$dummy [983]), .D (nx1963), .CLK (clk), .R (rst)) ;
    mux21_ni ix1964 (.Y (nx1963), .A0 (camera_module_cache_ram_155__0), .A1 (
             nx34216), .S0 (nx34328)) ;
    aoi22 ix28519 (.Y (nx28518), .A0 (camera_module_cache_ram_187__0), .A1 (
          nx36226), .B0 (camera_module_cache_ram_171__0), .B1 (nx36266)) ;
    dffr camera_module_cache_reg_ram_187__0 (.Q (camera_module_cache_ram_187__0)
         , .QB (\$dummy [984]), .D (nx1943), .CLK (clk), .R (rst)) ;
    mux21_ni ix1944 (.Y (nx1943), .A0 (camera_module_cache_ram_187__0), .A1 (
             nx34216), .S0 (nx34320)) ;
    dffr camera_module_cache_reg_ram_171__0 (.Q (camera_module_cache_ram_171__0)
         , .QB (\$dummy [985]), .D (nx1953), .CLK (clk), .R (rst)) ;
    mux21_ni ix1954 (.Y (nx1953), .A0 (camera_module_cache_ram_171__0), .A1 (
             nx34216), .S0 (nx34324)) ;
    aoi22 ix28527 (.Y (nx28526), .A0 (camera_module_cache_ram_203__0), .A1 (
          nx36306), .B0 (camera_module_cache_ram_219__0), .B1 (nx36346)) ;
    dffr camera_module_cache_reg_ram_203__0 (.Q (camera_module_cache_ram_203__0)
         , .QB (\$dummy [986]), .D (nx1933), .CLK (clk), .R (rst)) ;
    mux21_ni ix1934 (.Y (nx1933), .A0 (camera_module_cache_ram_203__0), .A1 (
             nx34216), .S0 (nx34316)) ;
    dffr camera_module_cache_reg_ram_219__0 (.Q (camera_module_cache_ram_219__0)
         , .QB (\$dummy [987]), .D (nx1923), .CLK (clk), .R (rst)) ;
    mux21_ni ix1924 (.Y (nx1923), .A0 (camera_module_cache_ram_219__0), .A1 (
             nx34218), .S0 (nx34312)) ;
    aoi22 ix28535 (.Y (nx28534), .A0 (camera_module_cache_ram_235__0), .A1 (
          nx36386), .B0 (camera_module_cache_ram_251__0), .B1 (nx36426)) ;
    dffr camera_module_cache_reg_ram_235__0 (.Q (camera_module_cache_ram_235__0)
         , .QB (\$dummy [988]), .D (nx1913), .CLK (clk), .R (rst)) ;
    mux21_ni ix1914 (.Y (nx1913), .A0 (camera_module_cache_ram_235__0), .A1 (
             nx34218), .S0 (nx34308)) ;
    dffr camera_module_cache_reg_ram_251__0 (.Q (camera_module_cache_ram_251__0)
         , .QB (\$dummy [989]), .D (nx1903), .CLK (clk), .R (rst)) ;
    mux21_ni ix1904 (.Y (nx1903), .A0 (camera_module_cache_ram_251__0), .A1 (
             nx34218), .S0 (nx34304)) ;
    nand04 ix2411 (.Y (nx2410), .A0 (nx28543), .A1 (nx28611), .A2 (nx28679), .A3 (
           nx28747)) ;
    oai21 ix28544 (.Y (nx28543), .A0 (nx2400), .A1 (nx2258), .B0 (nx36506)) ;
    nand04 ix2401 (.Y (nx2400), .A0 (nx28546), .A1 (nx28554), .A2 (nx28562), .A3 (
           nx28570)) ;
    aoi22 ix28547 (.Y (nx28546), .A0 (camera_module_cache_ram_12__0), .A1 (
          nx35826), .B0 (camera_module_cache_ram_28__0), .B1 (nx35866)) ;
    dffr camera_module_cache_reg_ram_12__0 (.Q (camera_module_cache_ram_12__0), 
         .QB (\$dummy [990]), .D (nx1893), .CLK (clk), .R (rst)) ;
    mux21_ni ix1894 (.Y (nx1893), .A0 (nx34218), .A1 (
             camera_module_cache_ram_12__0), .S0 (nx36496)) ;
    dffr camera_module_cache_reg_ram_28__0 (.Q (camera_module_cache_ram_28__0), 
         .QB (\$dummy [991]), .D (nx1883), .CLK (clk), .R (rst)) ;
    mux21_ni ix1884 (.Y (nx1883), .A0 (nx34218), .A1 (
             camera_module_cache_ram_28__0), .S0 (nx36510)) ;
    aoi22 ix28555 (.Y (nx28554), .A0 (camera_module_cache_ram_44__0), .A1 (
          nx35906), .B0 (camera_module_cache_ram_60__0), .B1 (nx35946)) ;
    dffr camera_module_cache_reg_ram_44__0 (.Q (camera_module_cache_ram_44__0), 
         .QB (\$dummy [992]), .D (nx1873), .CLK (clk), .R (rst)) ;
    mux21_ni ix1874 (.Y (nx1873), .A0 (nx34218), .A1 (
             camera_module_cache_ram_44__0), .S0 (nx36514)) ;
    dffr camera_module_cache_reg_ram_60__0 (.Q (camera_module_cache_ram_60__0), 
         .QB (\$dummy [993]), .D (nx1863), .CLK (clk), .R (rst)) ;
    mux21_ni ix1864 (.Y (nx1863), .A0 (nx34218), .A1 (
             camera_module_cache_ram_60__0), .S0 (nx36518)) ;
    aoi22 ix28563 (.Y (nx28562), .A0 (camera_module_cache_ram_76__0), .A1 (
          nx35986), .B0 (camera_module_cache_ram_92__0), .B1 (nx36026)) ;
    dffr camera_module_cache_reg_ram_76__0 (.Q (camera_module_cache_ram_76__0), 
         .QB (\$dummy [994]), .D (nx1853), .CLK (clk), .R (rst)) ;
    mux21_ni ix1854 (.Y (nx1853), .A0 (nx34220), .A1 (
             camera_module_cache_ram_76__0), .S0 (nx36522)) ;
    dffr camera_module_cache_reg_ram_92__0 (.Q (camera_module_cache_ram_92__0), 
         .QB (\$dummy [995]), .D (nx1843), .CLK (clk), .R (rst)) ;
    mux21_ni ix1844 (.Y (nx1843), .A0 (nx34220), .A1 (
             camera_module_cache_ram_92__0), .S0 (nx36526)) ;
    aoi22 ix28571 (.Y (nx28570), .A0 (camera_module_cache_ram_124__0), .A1 (
          nx36066), .B0 (camera_module_cache_ram_108__0), .B1 (nx36106)) ;
    dffr camera_module_cache_reg_ram_124__0 (.Q (camera_module_cache_ram_124__0)
         , .QB (\$dummy [996]), .D (nx1823), .CLK (clk), .R (rst)) ;
    mux21_ni ix1824 (.Y (nx1823), .A0 (nx34220), .A1 (
             camera_module_cache_ram_124__0), .S0 (nx36530)) ;
    dffr camera_module_cache_reg_ram_108__0 (.Q (camera_module_cache_ram_108__0)
         , .QB (\$dummy [997]), .D (nx1833), .CLK (clk), .R (rst)) ;
    mux21_ni ix1834 (.Y (nx1833), .A0 (nx34220), .A1 (
             camera_module_cache_ram_108__0), .S0 (nx36534)) ;
    nand04 ix2259 (.Y (nx2258), .A0 (nx28579), .A1 (nx28587), .A2 (nx28595), .A3 (
           nx28603)) ;
    aoi22 ix28580 (.Y (nx28579), .A0 (camera_module_cache_ram_140__0), .A1 (
          nx36146), .B0 (camera_module_cache_ram_156__0), .B1 (nx36186)) ;
    dffr camera_module_cache_reg_ram_140__0 (.Q (camera_module_cache_ram_140__0)
         , .QB (\$dummy [998]), .D (nx1813), .CLK (clk), .R (rst)) ;
    mux21_ni ix1814 (.Y (nx1813), .A0 (nx34220), .A1 (
             camera_module_cache_ram_140__0), .S0 (nx36538)) ;
    dffr camera_module_cache_reg_ram_156__0 (.Q (camera_module_cache_ram_156__0)
         , .QB (\$dummy [999]), .D (nx1803), .CLK (clk), .R (rst)) ;
    mux21_ni ix1804 (.Y (nx1803), .A0 (nx34220), .A1 (
             camera_module_cache_ram_156__0), .S0 (nx36542)) ;
    aoi22 ix28588 (.Y (nx28587), .A0 (camera_module_cache_ram_188__0), .A1 (
          nx36226), .B0 (camera_module_cache_ram_172__0), .B1 (nx36266)) ;
    dffr camera_module_cache_reg_ram_188__0 (.Q (camera_module_cache_ram_188__0)
         , .QB (\$dummy [1000]), .D (nx1783), .CLK (clk), .R (rst)) ;
    mux21_ni ix1784 (.Y (nx1783), .A0 (nx34220), .A1 (
             camera_module_cache_ram_188__0), .S0 (nx36546)) ;
    dffr camera_module_cache_reg_ram_172__0 (.Q (camera_module_cache_ram_172__0)
         , .QB (\$dummy [1001]), .D (nx1793), .CLK (clk), .R (rst)) ;
    mux21_ni ix1794 (.Y (nx1793), .A0 (nx34222), .A1 (
             camera_module_cache_ram_172__0), .S0 (nx36550)) ;
    aoi22 ix28596 (.Y (nx28595), .A0 (camera_module_cache_ram_204__0), .A1 (
          nx36306), .B0 (camera_module_cache_ram_220__0), .B1 (nx36346)) ;
    dffr camera_module_cache_reg_ram_204__0 (.Q (camera_module_cache_ram_204__0)
         , .QB (\$dummy [1002]), .D (nx1773), .CLK (clk), .R (rst)) ;
    mux21_ni ix1774 (.Y (nx1773), .A0 (nx34222), .A1 (
             camera_module_cache_ram_204__0), .S0 (nx36554)) ;
    dffr camera_module_cache_reg_ram_220__0 (.Q (camera_module_cache_ram_220__0)
         , .QB (\$dummy [1003]), .D (nx1763), .CLK (clk), .R (rst)) ;
    mux21_ni ix1764 (.Y (nx1763), .A0 (nx34222), .A1 (
             camera_module_cache_ram_220__0), .S0 (nx36558)) ;
    aoi22 ix28604 (.Y (nx28603), .A0 (camera_module_cache_ram_236__0), .A1 (
          nx36386), .B0 (camera_module_cache_ram_252__0), .B1 (nx36426)) ;
    dffr camera_module_cache_reg_ram_236__0 (.Q (camera_module_cache_ram_236__0)
         , .QB (\$dummy [1004]), .D (nx1753), .CLK (clk), .R (rst)) ;
    mux21_ni ix1754 (.Y (nx1753), .A0 (nx34222), .A1 (
             camera_module_cache_ram_236__0), .S0 (nx36562)) ;
    dffr camera_module_cache_reg_ram_252__0 (.Q (camera_module_cache_ram_252__0)
         , .QB (\$dummy [1005]), .D (nx1743), .CLK (clk), .R (rst)) ;
    mux21_ni ix1744 (.Y (nx1743), .A0 (nx34222), .A1 (
             camera_module_cache_ram_252__0), .S0 (nx36566)) ;
    oai21 ix28612 (.Y (nx28611), .A0 (nx2106), .A1 (nx1964), .B0 (nx36580)) ;
    nand04 ix2107 (.Y (nx2106), .A0 (nx28614), .A1 (nx28622), .A2 (nx28630), .A3 (
           nx28638)) ;
    aoi22 ix28615 (.Y (nx28614), .A0 (camera_module_cache_ram_13__0), .A1 (
          nx35826), .B0 (camera_module_cache_ram_29__0), .B1 (nx35866)) ;
    dffr camera_module_cache_reg_ram_13__0 (.Q (camera_module_cache_ram_13__0), 
         .QB (\$dummy [1006]), .D (nx1733), .CLK (clk), .R (rst)) ;
    mux21_ni ix1734 (.Y (nx1733), .A0 (nx34222), .A1 (
             camera_module_cache_ram_13__0), .S0 (nx36570)) ;
    dffr camera_module_cache_reg_ram_29__0 (.Q (camera_module_cache_ram_29__0), 
         .QB (\$dummy [1007]), .D (nx1723), .CLK (clk), .R (rst)) ;
    mux21_ni ix1724 (.Y (nx1723), .A0 (nx34222), .A1 (
             camera_module_cache_ram_29__0), .S0 (nx36584)) ;
    aoi22 ix28623 (.Y (nx28622), .A0 (camera_module_cache_ram_45__0), .A1 (
          nx35906), .B0 (camera_module_cache_ram_61__0), .B1 (nx35946)) ;
    dffr camera_module_cache_reg_ram_45__0 (.Q (camera_module_cache_ram_45__0), 
         .QB (\$dummy [1008]), .D (nx1713), .CLK (clk), .R (rst)) ;
    mux21_ni ix1714 (.Y (nx1713), .A0 (nx34224), .A1 (
             camera_module_cache_ram_45__0), .S0 (nx36588)) ;
    dffr camera_module_cache_reg_ram_61__0 (.Q (camera_module_cache_ram_61__0), 
         .QB (\$dummy [1009]), .D (nx1703), .CLK (clk), .R (rst)) ;
    mux21_ni ix1704 (.Y (nx1703), .A0 (nx34224), .A1 (
             camera_module_cache_ram_61__0), .S0 (nx36592)) ;
    aoi22 ix28631 (.Y (nx28630), .A0 (camera_module_cache_ram_77__0), .A1 (
          nx35986), .B0 (camera_module_cache_ram_93__0), .B1 (nx36026)) ;
    dffr camera_module_cache_reg_ram_77__0 (.Q (camera_module_cache_ram_77__0), 
         .QB (\$dummy [1010]), .D (nx1693), .CLK (clk), .R (rst)) ;
    mux21_ni ix1694 (.Y (nx1693), .A0 (nx34224), .A1 (
             camera_module_cache_ram_77__0), .S0 (nx36596)) ;
    dffr camera_module_cache_reg_ram_93__0 (.Q (camera_module_cache_ram_93__0), 
         .QB (\$dummy [1011]), .D (nx1683), .CLK (clk), .R (rst)) ;
    mux21_ni ix1684 (.Y (nx1683), .A0 (nx34224), .A1 (
             camera_module_cache_ram_93__0), .S0 (nx36600)) ;
    aoi22 ix28639 (.Y (nx28638), .A0 (camera_module_cache_ram_125__0), .A1 (
          nx36066), .B0 (camera_module_cache_ram_109__0), .B1 (nx36106)) ;
    dffr camera_module_cache_reg_ram_125__0 (.Q (camera_module_cache_ram_125__0)
         , .QB (\$dummy [1012]), .D (nx1663), .CLK (clk), .R (rst)) ;
    mux21_ni ix1664 (.Y (nx1663), .A0 (nx34224), .A1 (
             camera_module_cache_ram_125__0), .S0 (nx36604)) ;
    dffr camera_module_cache_reg_ram_109__0 (.Q (camera_module_cache_ram_109__0)
         , .QB (\$dummy [1013]), .D (nx1673), .CLK (clk), .R (rst)) ;
    mux21_ni ix1674 (.Y (nx1673), .A0 (nx34224), .A1 (
             camera_module_cache_ram_109__0), .S0 (nx36608)) ;
    nand04 ix1965 (.Y (nx1964), .A0 (nx28647), .A1 (nx28655), .A2 (nx28663), .A3 (
           nx28671)) ;
    aoi22 ix28648 (.Y (nx28647), .A0 (camera_module_cache_ram_141__0), .A1 (
          nx36146), .B0 (camera_module_cache_ram_157__0), .B1 (nx36186)) ;
    dffr camera_module_cache_reg_ram_141__0 (.Q (camera_module_cache_ram_141__0)
         , .QB (\$dummy [1014]), .D (nx1653), .CLK (clk), .R (rst)) ;
    mux21_ni ix1654 (.Y (nx1653), .A0 (nx34224), .A1 (
             camera_module_cache_ram_141__0), .S0 (nx36612)) ;
    dffr camera_module_cache_reg_ram_157__0 (.Q (camera_module_cache_ram_157__0)
         , .QB (\$dummy [1015]), .D (nx1643), .CLK (clk), .R (rst)) ;
    mux21_ni ix1644 (.Y (nx1643), .A0 (nx34226), .A1 (
             camera_module_cache_ram_157__0), .S0 (nx36616)) ;
    aoi22 ix28656 (.Y (nx28655), .A0 (camera_module_cache_ram_189__0), .A1 (
          nx36226), .B0 (camera_module_cache_ram_173__0), .B1 (nx36266)) ;
    dffr camera_module_cache_reg_ram_189__0 (.Q (camera_module_cache_ram_189__0)
         , .QB (\$dummy [1016]), .D (nx1623), .CLK (clk), .R (rst)) ;
    mux21_ni ix1624 (.Y (nx1623), .A0 (nx34226), .A1 (
             camera_module_cache_ram_189__0), .S0 (nx36620)) ;
    dffr camera_module_cache_reg_ram_173__0 (.Q (camera_module_cache_ram_173__0)
         , .QB (\$dummy [1017]), .D (nx1633), .CLK (clk), .R (rst)) ;
    mux21_ni ix1634 (.Y (nx1633), .A0 (nx34226), .A1 (
             camera_module_cache_ram_173__0), .S0 (nx36624)) ;
    aoi22 ix28664 (.Y (nx28663), .A0 (camera_module_cache_ram_205__0), .A1 (
          nx36306), .B0 (camera_module_cache_ram_221__0), .B1 (nx36346)) ;
    dffr camera_module_cache_reg_ram_205__0 (.Q (camera_module_cache_ram_205__0)
         , .QB (\$dummy [1018]), .D (nx1613), .CLK (clk), .R (rst)) ;
    mux21_ni ix1614 (.Y (nx1613), .A0 (nx34226), .A1 (
             camera_module_cache_ram_205__0), .S0 (nx36628)) ;
    dffr camera_module_cache_reg_ram_221__0 (.Q (camera_module_cache_ram_221__0)
         , .QB (\$dummy [1019]), .D (nx1603), .CLK (clk), .R (rst)) ;
    mux21_ni ix1604 (.Y (nx1603), .A0 (nx34226), .A1 (
             camera_module_cache_ram_221__0), .S0 (nx36632)) ;
    aoi22 ix28672 (.Y (nx28671), .A0 (camera_module_cache_ram_237__0), .A1 (
          nx36386), .B0 (camera_module_cache_ram_253__0), .B1 (nx36426)) ;
    dffr camera_module_cache_reg_ram_237__0 (.Q (camera_module_cache_ram_237__0)
         , .QB (\$dummy [1020]), .D (nx1593), .CLK (clk), .R (rst)) ;
    mux21_ni ix1594 (.Y (nx1593), .A0 (nx34226), .A1 (
             camera_module_cache_ram_237__0), .S0 (nx36636)) ;
    dffr camera_module_cache_reg_ram_253__0 (.Q (camera_module_cache_ram_253__0)
         , .QB (\$dummy [1021]), .D (nx1583), .CLK (clk), .R (rst)) ;
    mux21_ni ix1584 (.Y (nx1583), .A0 (nx34226), .A1 (
             camera_module_cache_ram_253__0), .S0 (nx36640)) ;
    oai21 ix28680 (.Y (nx28679), .A0 (nx1808), .A1 (nx1666), .B0 (nx36654)) ;
    nand04 ix1809 (.Y (nx1808), .A0 (nx28682), .A1 (nx28690), .A2 (nx28698), .A3 (
           nx28706)) ;
    aoi22 ix28683 (.Y (nx28682), .A0 (camera_module_cache_ram_14__0), .A1 (
          nx35826), .B0 (camera_module_cache_ram_30__0), .B1 (nx35866)) ;
    dffr camera_module_cache_reg_ram_14__0 (.Q (camera_module_cache_ram_14__0), 
         .QB (\$dummy [1022]), .D (nx1573), .CLK (clk), .R (rst)) ;
    mux21_ni ix1574 (.Y (nx1573), .A0 (nx34228), .A1 (
             camera_module_cache_ram_14__0), .S0 (nx36644)) ;
    dffr camera_module_cache_reg_ram_30__0 (.Q (camera_module_cache_ram_30__0), 
         .QB (\$dummy [1023]), .D (nx1563), .CLK (clk), .R (rst)) ;
    mux21_ni ix1564 (.Y (nx1563), .A0 (nx34228), .A1 (
             camera_module_cache_ram_30__0), .S0 (nx36658)) ;
    aoi22 ix28691 (.Y (nx28690), .A0 (camera_module_cache_ram_46__0), .A1 (
          nx35906), .B0 (camera_module_cache_ram_62__0), .B1 (nx35946)) ;
    dffr camera_module_cache_reg_ram_46__0 (.Q (camera_module_cache_ram_46__0), 
         .QB (\$dummy [1024]), .D (nx1553), .CLK (clk), .R (rst)) ;
    mux21_ni ix1554 (.Y (nx1553), .A0 (nx34228), .A1 (
             camera_module_cache_ram_46__0), .S0 (nx36662)) ;
    dffr camera_module_cache_reg_ram_62__0 (.Q (camera_module_cache_ram_62__0), 
         .QB (\$dummy [1025]), .D (nx1543), .CLK (clk), .R (rst)) ;
    mux21_ni ix1544 (.Y (nx1543), .A0 (nx34228), .A1 (
             camera_module_cache_ram_62__0), .S0 (nx36666)) ;
    aoi22 ix28699 (.Y (nx28698), .A0 (camera_module_cache_ram_78__0), .A1 (
          nx35986), .B0 (camera_module_cache_ram_94__0), .B1 (nx36026)) ;
    dffr camera_module_cache_reg_ram_78__0 (.Q (camera_module_cache_ram_78__0), 
         .QB (\$dummy [1026]), .D (nx1533), .CLK (clk), .R (rst)) ;
    mux21_ni ix1534 (.Y (nx1533), .A0 (nx34228), .A1 (
             camera_module_cache_ram_78__0), .S0 (nx36670)) ;
    dffr camera_module_cache_reg_ram_94__0 (.Q (camera_module_cache_ram_94__0), 
         .QB (\$dummy [1027]), .D (nx1523), .CLK (clk), .R (rst)) ;
    mux21_ni ix1524 (.Y (nx1523), .A0 (nx34228), .A1 (
             camera_module_cache_ram_94__0), .S0 (nx36674)) ;
    aoi22 ix28707 (.Y (nx28706), .A0 (camera_module_cache_ram_126__0), .A1 (
          nx36066), .B0 (camera_module_cache_ram_110__0), .B1 (nx36106)) ;
    dffr camera_module_cache_reg_ram_126__0 (.Q (camera_module_cache_ram_126__0)
         , .QB (\$dummy [1028]), .D (nx1503), .CLK (clk), .R (rst)) ;
    mux21_ni ix1504 (.Y (nx1503), .A0 (nx34228), .A1 (
             camera_module_cache_ram_126__0), .S0 (nx36678)) ;
    dffr camera_module_cache_reg_ram_110__0 (.Q (camera_module_cache_ram_110__0)
         , .QB (\$dummy [1029]), .D (nx1513), .CLK (clk), .R (rst)) ;
    mux21_ni ix1514 (.Y (nx1513), .A0 (nx34230), .A1 (
             camera_module_cache_ram_110__0), .S0 (nx36682)) ;
    nand04 ix1667 (.Y (nx1666), .A0 (nx28715), .A1 (nx28723), .A2 (nx28731), .A3 (
           nx28739)) ;
    aoi22 ix28716 (.Y (nx28715), .A0 (camera_module_cache_ram_142__0), .A1 (
          nx36146), .B0 (camera_module_cache_ram_158__0), .B1 (nx36186)) ;
    dffr camera_module_cache_reg_ram_142__0 (.Q (camera_module_cache_ram_142__0)
         , .QB (\$dummy [1030]), .D (nx1493), .CLK (clk), .R (rst)) ;
    mux21_ni ix1494 (.Y (nx1493), .A0 (nx34230), .A1 (
             camera_module_cache_ram_142__0), .S0 (nx36686)) ;
    dffr camera_module_cache_reg_ram_158__0 (.Q (camera_module_cache_ram_158__0)
         , .QB (\$dummy [1031]), .D (nx1483), .CLK (clk), .R (rst)) ;
    mux21_ni ix1484 (.Y (nx1483), .A0 (nx34230), .A1 (
             camera_module_cache_ram_158__0), .S0 (nx36690)) ;
    aoi22 ix28724 (.Y (nx28723), .A0 (camera_module_cache_ram_190__0), .A1 (
          nx36226), .B0 (camera_module_cache_ram_174__0), .B1 (nx36266)) ;
    dffr camera_module_cache_reg_ram_190__0 (.Q (camera_module_cache_ram_190__0)
         , .QB (\$dummy [1032]), .D (nx1463), .CLK (clk), .R (rst)) ;
    mux21_ni ix1464 (.Y (nx1463), .A0 (nx34230), .A1 (
             camera_module_cache_ram_190__0), .S0 (nx36694)) ;
    dffr camera_module_cache_reg_ram_174__0 (.Q (camera_module_cache_ram_174__0)
         , .QB (\$dummy [1033]), .D (nx1473), .CLK (clk), .R (rst)) ;
    mux21_ni ix1474 (.Y (nx1473), .A0 (nx34230), .A1 (
             camera_module_cache_ram_174__0), .S0 (nx36698)) ;
    aoi22 ix28732 (.Y (nx28731), .A0 (camera_module_cache_ram_206__0), .A1 (
          nx36306), .B0 (camera_module_cache_ram_222__0), .B1 (nx36346)) ;
    dffr camera_module_cache_reg_ram_206__0 (.Q (camera_module_cache_ram_206__0)
         , .QB (\$dummy [1034]), .D (nx1453), .CLK (clk), .R (rst)) ;
    mux21_ni ix1454 (.Y (nx1453), .A0 (nx34230), .A1 (
             camera_module_cache_ram_206__0), .S0 (nx36702)) ;
    dffr camera_module_cache_reg_ram_222__0 (.Q (camera_module_cache_ram_222__0)
         , .QB (\$dummy [1035]), .D (nx1443), .CLK (clk), .R (rst)) ;
    mux21_ni ix1444 (.Y (nx1443), .A0 (nx34230), .A1 (
             camera_module_cache_ram_222__0), .S0 (nx36706)) ;
    aoi22 ix28740 (.Y (nx28739), .A0 (camera_module_cache_ram_238__0), .A1 (
          nx36386), .B0 (camera_module_cache_ram_254__0), .B1 (nx36426)) ;
    dffr camera_module_cache_reg_ram_238__0 (.Q (camera_module_cache_ram_238__0)
         , .QB (\$dummy [1036]), .D (nx1433), .CLK (clk), .R (rst)) ;
    mux21_ni ix1434 (.Y (nx1433), .A0 (nx34232), .A1 (
             camera_module_cache_ram_238__0), .S0 (nx36710)) ;
    dffr camera_module_cache_reg_ram_254__0 (.Q (camera_module_cache_ram_254__0)
         , .QB (\$dummy [1037]), .D (nx1423), .CLK (clk), .R (rst)) ;
    mux21_ni ix1424 (.Y (nx1423), .A0 (nx34232), .A1 (
             camera_module_cache_ram_254__0), .S0 (nx36714)) ;
    oai21 ix28748 (.Y (nx28747), .A0 (nx1512), .A1 (nx1348), .B0 (nx36728)) ;
    nand04 ix1513 (.Y (nx1512), .A0 (nx28750), .A1 (nx28758), .A2 (nx28766), .A3 (
           nx28774)) ;
    aoi22 ix28751 (.Y (nx28750), .A0 (camera_module_cache_ram_15__0), .A1 (
          nx35826), .B0 (camera_module_cache_ram_31__0), .B1 (nx35866)) ;
    dffr camera_module_cache_reg_ram_15__0 (.Q (camera_module_cache_ram_15__0), 
         .QB (\$dummy [1038]), .D (nx1413), .CLK (clk), .R (rst)) ;
    mux21_ni ix1414 (.Y (nx1413), .A0 (nx34232), .A1 (
             camera_module_cache_ram_15__0), .S0 (nx36718)) ;
    dffr camera_module_cache_reg_ram_31__0 (.Q (camera_module_cache_ram_31__0), 
         .QB (\$dummy [1039]), .D (nx1403), .CLK (clk), .R (rst)) ;
    mux21_ni ix1404 (.Y (nx1403), .A0 (nx34232), .A1 (
             camera_module_cache_ram_31__0), .S0 (nx36732)) ;
    aoi22 ix28759 (.Y (nx28758), .A0 (camera_module_cache_ram_47__0), .A1 (
          nx35906), .B0 (camera_module_cache_ram_63__0), .B1 (nx35946)) ;
    dffr camera_module_cache_reg_ram_47__0 (.Q (camera_module_cache_ram_47__0), 
         .QB (\$dummy [1040]), .D (nx1393), .CLK (clk), .R (rst)) ;
    mux21_ni ix1394 (.Y (nx1393), .A0 (nx34232), .A1 (
             camera_module_cache_ram_47__0), .S0 (nx36736)) ;
    dffr camera_module_cache_reg_ram_63__0 (.Q (camera_module_cache_ram_63__0), 
         .QB (\$dummy [1041]), .D (nx1383), .CLK (clk), .R (rst)) ;
    mux21_ni ix1384 (.Y (nx1383), .A0 (nx34232), .A1 (
             camera_module_cache_ram_63__0), .S0 (nx36740)) ;
    aoi22 ix28767 (.Y (nx28766), .A0 (camera_module_cache_ram_79__0), .A1 (
          nx35986), .B0 (camera_module_cache_ram_95__0), .B1 (nx36026)) ;
    dffr camera_module_cache_reg_ram_79__0 (.Q (camera_module_cache_ram_79__0), 
         .QB (\$dummy [1042]), .D (nx1373), .CLK (clk), .R (rst)) ;
    mux21_ni ix1374 (.Y (nx1373), .A0 (nx34232), .A1 (
             camera_module_cache_ram_79__0), .S0 (nx36744)) ;
    dffr camera_module_cache_reg_ram_95__0 (.Q (camera_module_cache_ram_95__0), 
         .QB (\$dummy [1043]), .D (nx1363), .CLK (clk), .R (rst)) ;
    mux21_ni ix1364 (.Y (nx1363), .A0 (nx34234), .A1 (
             camera_module_cache_ram_95__0), .S0 (nx36748)) ;
    aoi22 ix28775 (.Y (nx28774), .A0 (camera_module_cache_ram_127__0), .A1 (
          nx36066), .B0 (camera_module_cache_ram_111__0), .B1 (nx36106)) ;
    dffr camera_module_cache_reg_ram_127__0 (.Q (camera_module_cache_ram_127__0)
         , .QB (\$dummy [1044]), .D (nx1343), .CLK (clk), .R (rst)) ;
    mux21_ni ix1344 (.Y (nx1343), .A0 (nx34234), .A1 (
             camera_module_cache_ram_127__0), .S0 (nx36752)) ;
    dffr camera_module_cache_reg_ram_111__0 (.Q (camera_module_cache_ram_111__0)
         , .QB (\$dummy [1045]), .D (nx1353), .CLK (clk), .R (rst)) ;
    mux21_ni ix1354 (.Y (nx1353), .A0 (nx34234), .A1 (
             camera_module_cache_ram_111__0), .S0 (nx36756)) ;
    nand04 ix1349 (.Y (nx1348), .A0 (nx28783), .A1 (nx28791), .A2 (nx28799), .A3 (
           nx28807)) ;
    aoi22 ix28784 (.Y (nx28783), .A0 (camera_module_cache_ram_143__0), .A1 (
          nx36146), .B0 (camera_module_cache_ram_159__0), .B1 (nx36186)) ;
    dffr camera_module_cache_reg_ram_143__0 (.Q (camera_module_cache_ram_143__0)
         , .QB (\$dummy [1046]), .D (nx1333), .CLK (clk), .R (rst)) ;
    mux21_ni ix1334 (.Y (nx1333), .A0 (nx34234), .A1 (
             camera_module_cache_ram_143__0), .S0 (nx36760)) ;
    dffr camera_module_cache_reg_ram_159__0 (.Q (camera_module_cache_ram_159__0)
         , .QB (\$dummy [1047]), .D (nx1323), .CLK (clk), .R (rst)) ;
    mux21_ni ix1324 (.Y (nx1323), .A0 (nx34234), .A1 (
             camera_module_cache_ram_159__0), .S0 (nx36764)) ;
    aoi22 ix28792 (.Y (nx28791), .A0 (camera_module_cache_ram_191__0), .A1 (
          nx36226), .B0 (camera_module_cache_ram_175__0), .B1 (nx36266)) ;
    dffr camera_module_cache_reg_ram_191__0 (.Q (camera_module_cache_ram_191__0)
         , .QB (\$dummy [1048]), .D (nx1303), .CLK (clk), .R (rst)) ;
    mux21_ni ix1304 (.Y (nx1303), .A0 (nx34234), .A1 (
             camera_module_cache_ram_191__0), .S0 (nx36768)) ;
    dffr camera_module_cache_reg_ram_175__0 (.Q (camera_module_cache_ram_175__0)
         , .QB (\$dummy [1049]), .D (nx1313), .CLK (clk), .R (rst)) ;
    mux21_ni ix1314 (.Y (nx1313), .A0 (nx34234), .A1 (
             camera_module_cache_ram_175__0), .S0 (nx36772)) ;
    aoi22 ix28800 (.Y (nx28799), .A0 (camera_module_cache_ram_207__0), .A1 (
          nx36306), .B0 (camera_module_cache_ram_223__0), .B1 (nx36346)) ;
    dffr camera_module_cache_reg_ram_207__0 (.Q (camera_module_cache_ram_207__0)
         , .QB (\$dummy [1050]), .D (nx1293), .CLK (clk), .R (rst)) ;
    mux21_ni ix1294 (.Y (nx1293), .A0 (nx34236), .A1 (
             camera_module_cache_ram_207__0), .S0 (nx36776)) ;
    dffr camera_module_cache_reg_ram_223__0 (.Q (camera_module_cache_ram_223__0)
         , .QB (\$dummy [1051]), .D (nx1283), .CLK (clk), .R (rst)) ;
    mux21_ni ix1284 (.Y (nx1283), .A0 (nx34236), .A1 (
             camera_module_cache_ram_223__0), .S0 (nx36780)) ;
    aoi22 ix28808 (.Y (nx28807), .A0 (camera_module_cache_ram_239__0), .A1 (
          nx36386), .B0 (camera_module_cache_ram_255__0), .B1 (nx36426)) ;
    dffr camera_module_cache_reg_ram_239__0 (.Q (camera_module_cache_ram_239__0)
         , .QB (\$dummy [1052]), .D (nx1273), .CLK (clk), .R (rst)) ;
    mux21_ni ix1274 (.Y (nx1273), .A0 (nx34236), .A1 (
             camera_module_cache_ram_239__0), .S0 (nx36784)) ;
    dffr camera_module_cache_reg_ram_255__0 (.Q (camera_module_cache_ram_255__0)
         , .QB (\$dummy [1053]), .D (nx1263), .CLK (clk), .R (rst)) ;
    mux21_ni ix1264 (.Y (nx1263), .A0 (nx34236), .A1 (
             camera_module_cache_ram_255__0), .S0 (nx36788)) ;
    dff camera_module_algo_module_pixel_reg_reg_q_1 (.Q (
        camera_module_algo_module_pixel_value_1), .QB (nx29956), .D (nx6393), .CLK (
        clk)) ;
    mux21_ni ix6394 (.Y (nx6393), .A0 (nx8738), .A1 (
             camera_module_algo_module_pixel_value_1), .S0 (nx37152)) ;
    mux21_ni ix28823 (.Y (nx28822), .A0 (nx28824), .A1 (nx35676), .S0 (nx36792)
             ) ;
    nor04 ix28825 (.Y (nx28824), .A0 (nx8718), .A1 (nx8064), .A2 (nx7408), .A3 (
          nx6754)) ;
    nand04 ix8719 (.Y (nx8718), .A0 (nx28827), .A1 (nx28933), .A2 (nx29001), .A3 (
           nx29069)) ;
    oai21 ix28828 (.Y (nx28827), .A0 (nx8708), .A1 (nx8630), .B0 (nx36448)) ;
    nand04 ix8709 (.Y (nx8708), .A0 (nx28830), .A1 (nx28876), .A2 (nx28884), .A3 (
           nx28892)) ;
    aoi22 ix28831 (.Y (nx28830), .A0 (camera_module_cache_ram_0__1), .A1 (
          nx35826), .B0 (camera_module_cache_ram_16__1), .B1 (nx35866)) ;
    dffr camera_module_cache_reg_ram_0__1 (.Q (camera_module_cache_ram_0__1), .QB (
         \$dummy [1054]), .D (nx6383), .CLK (clk), .R (rst)) ;
    mux21_ni ix6384 (.Y (nx6383), .A0 (camera_module_cache_ram_0__1), .A1 (
             nx35140), .S0 (nx35134)) ;
    oai221 ix6101 (.Y (nx6100), .A0 (nx34074), .A1 (nx28835), .B0 (nx28851), .B1 (
           nx35712), .C0 (nx28854)) ;
    tri01 nvm_module_tri_dataout_121 (.Y (nvm_data_121), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_113 (.Y (nvm_data_113), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_105 (.Y (nvm_data_105), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_97 (.Y (nvm_data_97), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_89 (.Y (nvm_data_89), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_81 (.Y (nvm_data_81), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_73 (.Y (nvm_data_73), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_65 (.Y (nvm_data_65), .A (nx22549), .E (
          nvm_module_GND0)) ;
    inv01 ix28852 (.Y (nx28851), .A (nvm_data_1)) ;
    tri01 nvm_module_tri_dataout_1 (.Y (nvm_data_1), .A (nx22549), .E (
          nvm_module_GND0)) ;
    nand02 ix28855 (.Y (nx28854), .A0 (nx34074), .A1 (nx6034)) ;
    tri01 nvm_module_tri_dataout_57 (.Y (nvm_data_57), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_49 (.Y (nvm_data_49), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_41 (.Y (nvm_data_41), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_33 (.Y (nvm_data_33), .A (nx22549), .E (
          nvm_module_GND0)) ;
    oai22 ix6003 (.Y (nx6002), .A0 (nx34104), .A1 (nx28865), .B0 (nx34090), .B1 (
          nx28869)) ;
    tri01 nvm_module_tri_dataout_25 (.Y (nvm_data_25), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_17 (.Y (nvm_data_17), .A (nx22549), .E (
          nvm_module_GND0)) ;
    nand02 ix28870 (.Y (nx28869), .A0 (nvm_data_9), .A1 (nx34106)) ;
    tri01 nvm_module_tri_dataout_9 (.Y (nvm_data_9), .A (nx22549), .E (
          nvm_module_GND0)) ;
    dffr camera_module_cache_reg_ram_16__1 (.Q (camera_module_cache_ram_16__1), 
         .QB (\$dummy [1055]), .D (nx6373), .CLK (clk), .R (rst)) ;
    mux21_ni ix6374 (.Y (nx6373), .A0 (camera_module_cache_ram_16__1), .A1 (
             nx35140), .S0 (nx35130)) ;
    aoi22 ix28877 (.Y (nx28876), .A0 (camera_module_cache_ram_32__1), .A1 (
          nx35906), .B0 (camera_module_cache_ram_48__1), .B1 (nx35946)) ;
    dffr camera_module_cache_reg_ram_32__1 (.Q (camera_module_cache_ram_32__1), 
         .QB (\$dummy [1056]), .D (nx6363), .CLK (clk), .R (rst)) ;
    mux21_ni ix6364 (.Y (nx6363), .A0 (camera_module_cache_ram_32__1), .A1 (
             nx35140), .S0 (nx35126)) ;
    dffr camera_module_cache_reg_ram_48__1 (.Q (camera_module_cache_ram_48__1), 
         .QB (\$dummy [1057]), .D (nx6353), .CLK (clk), .R (rst)) ;
    mux21_ni ix6354 (.Y (nx6353), .A0 (camera_module_cache_ram_48__1), .A1 (
             nx35140), .S0 (nx35122)) ;
    aoi22 ix28885 (.Y (nx28884), .A0 (camera_module_cache_ram_64__1), .A1 (
          nx35986), .B0 (camera_module_cache_ram_80__1), .B1 (nx36026)) ;
    dffr camera_module_cache_reg_ram_64__1 (.Q (camera_module_cache_ram_64__1), 
         .QB (\$dummy [1058]), .D (nx6343), .CLK (clk), .R (rst)) ;
    mux21_ni ix6344 (.Y (nx6343), .A0 (camera_module_cache_ram_64__1), .A1 (
             nx35140), .S0 (nx35118)) ;
    dffr camera_module_cache_reg_ram_80__1 (.Q (camera_module_cache_ram_80__1), 
         .QB (\$dummy [1059]), .D (nx6333), .CLK (clk), .R (rst)) ;
    mux21_ni ix6334 (.Y (nx6333), .A0 (camera_module_cache_ram_80__1), .A1 (
             nx35140), .S0 (nx35114)) ;
    aoi22 ix28893 (.Y (nx28892), .A0 (camera_module_cache_ram_112__1), .A1 (
          nx36066), .B0 (camera_module_cache_ram_96__1), .B1 (nx36106)) ;
    dffr camera_module_cache_reg_ram_112__1 (.Q (camera_module_cache_ram_112__1)
         , .QB (\$dummy [1060]), .D (nx6313), .CLK (clk), .R (rst)) ;
    mux21_ni ix6314 (.Y (nx6313), .A0 (camera_module_cache_ram_112__1), .A1 (
             nx35140), .S0 (nx35106)) ;
    dffr camera_module_cache_reg_ram_96__1 (.Q (camera_module_cache_ram_96__1), 
         .QB (\$dummy [1061]), .D (nx6323), .CLK (clk), .R (rst)) ;
    mux21_ni ix6324 (.Y (nx6323), .A0 (camera_module_cache_ram_96__1), .A1 (
             nx35142), .S0 (nx35110)) ;
    nand04 ix8631 (.Y (nx8630), .A0 (nx28901), .A1 (nx28909), .A2 (nx28917), .A3 (
           nx28925)) ;
    aoi22 ix28902 (.Y (nx28901), .A0 (camera_module_cache_ram_128__1), .A1 (
          nx36146), .B0 (camera_module_cache_ram_144__1), .B1 (nx36186)) ;
    dffr camera_module_cache_reg_ram_128__1 (.Q (camera_module_cache_ram_128__1)
         , .QB (\$dummy [1062]), .D (nx6303), .CLK (clk), .R (rst)) ;
    mux21_ni ix6304 (.Y (nx6303), .A0 (camera_module_cache_ram_128__1), .A1 (
             nx35142), .S0 (nx35102)) ;
    dffr camera_module_cache_reg_ram_144__1 (.Q (camera_module_cache_ram_144__1)
         , .QB (\$dummy [1063]), .D (nx6293), .CLK (clk), .R (rst)) ;
    mux21_ni ix6294 (.Y (nx6293), .A0 (camera_module_cache_ram_144__1), .A1 (
             nx35142), .S0 (nx35098)) ;
    aoi22 ix28910 (.Y (nx28909), .A0 (camera_module_cache_ram_176__1), .A1 (
          nx36226), .B0 (camera_module_cache_ram_160__1), .B1 (nx36266)) ;
    dffr camera_module_cache_reg_ram_176__1 (.Q (camera_module_cache_ram_176__1)
         , .QB (\$dummy [1064]), .D (nx6273), .CLK (clk), .R (rst)) ;
    mux21_ni ix6274 (.Y (nx6273), .A0 (camera_module_cache_ram_176__1), .A1 (
             nx35142), .S0 (nx35090)) ;
    dffr camera_module_cache_reg_ram_160__1 (.Q (camera_module_cache_ram_160__1)
         , .QB (\$dummy [1065]), .D (nx6283), .CLK (clk), .R (rst)) ;
    mux21_ni ix6284 (.Y (nx6283), .A0 (camera_module_cache_ram_160__1), .A1 (
             nx35142), .S0 (nx35094)) ;
    aoi22 ix28918 (.Y (nx28917), .A0 (camera_module_cache_ram_192__1), .A1 (
          nx36306), .B0 (camera_module_cache_ram_208__1), .B1 (nx36346)) ;
    dffr camera_module_cache_reg_ram_192__1 (.Q (camera_module_cache_ram_192__1)
         , .QB (\$dummy [1066]), .D (nx6263), .CLK (clk), .R (rst)) ;
    mux21_ni ix6264 (.Y (nx6263), .A0 (camera_module_cache_ram_192__1), .A1 (
             nx35142), .S0 (nx35086)) ;
    dffr camera_module_cache_reg_ram_208__1 (.Q (camera_module_cache_ram_208__1)
         , .QB (\$dummy [1067]), .D (nx6253), .CLK (clk), .R (rst)) ;
    mux21_ni ix6254 (.Y (nx6253), .A0 (camera_module_cache_ram_208__1), .A1 (
             nx35142), .S0 (nx35082)) ;
    aoi22 ix28926 (.Y (nx28925), .A0 (camera_module_cache_ram_224__1), .A1 (
          nx36386), .B0 (camera_module_cache_ram_240__1), .B1 (nx36426)) ;
    dffr camera_module_cache_reg_ram_224__1 (.Q (camera_module_cache_ram_224__1)
         , .QB (\$dummy [1068]), .D (nx6243), .CLK (clk), .R (rst)) ;
    mux21_ni ix6244 (.Y (nx6243), .A0 (camera_module_cache_ram_224__1), .A1 (
             nx35144), .S0 (nx35078)) ;
    dffr camera_module_cache_reg_ram_240__1 (.Q (camera_module_cache_ram_240__1)
         , .QB (\$dummy [1069]), .D (nx6233), .CLK (clk), .R (rst)) ;
    mux21_ni ix6234 (.Y (nx6233), .A0 (camera_module_cache_ram_240__1), .A1 (
             nx35144), .S0 (nx35074)) ;
    oai21 ix28934 (.Y (nx28933), .A0 (nx8546), .A1 (nx8468), .B0 (nx36452)) ;
    nand04 ix8547 (.Y (nx8546), .A0 (nx28936), .A1 (nx28944), .A2 (nx28952), .A3 (
           nx28960)) ;
    aoi22 ix28937 (.Y (nx28936), .A0 (camera_module_cache_ram_1__1), .A1 (
          nx35826), .B0 (camera_module_cache_ram_17__1), .B1 (nx35866)) ;
    dffr camera_module_cache_reg_ram_1__1 (.Q (camera_module_cache_ram_1__1), .QB (
         \$dummy [1070]), .D (nx6223), .CLK (clk), .R (rst)) ;
    mux21_ni ix6224 (.Y (nx6223), .A0 (camera_module_cache_ram_1__1), .A1 (
             nx35144), .S0 (nx35064)) ;
    dffr camera_module_cache_reg_ram_17__1 (.Q (camera_module_cache_ram_17__1), 
         .QB (\$dummy [1071]), .D (nx6213), .CLK (clk), .R (rst)) ;
    mux21_ni ix6214 (.Y (nx6213), .A0 (camera_module_cache_ram_17__1), .A1 (
             nx35144), .S0 (nx35060)) ;
    aoi22 ix28945 (.Y (nx28944), .A0 (camera_module_cache_ram_33__1), .A1 (
          nx35906), .B0 (camera_module_cache_ram_49__1), .B1 (nx35946)) ;
    dffr camera_module_cache_reg_ram_33__1 (.Q (camera_module_cache_ram_33__1), 
         .QB (\$dummy [1072]), .D (nx6203), .CLK (clk), .R (rst)) ;
    mux21_ni ix6204 (.Y (nx6203), .A0 (camera_module_cache_ram_33__1), .A1 (
             nx35144), .S0 (nx35056)) ;
    dffr camera_module_cache_reg_ram_49__1 (.Q (camera_module_cache_ram_49__1), 
         .QB (\$dummy [1073]), .D (nx6193), .CLK (clk), .R (rst)) ;
    mux21_ni ix6194 (.Y (nx6193), .A0 (camera_module_cache_ram_49__1), .A1 (
             nx35144), .S0 (nx35052)) ;
    aoi22 ix28953 (.Y (nx28952), .A0 (camera_module_cache_ram_65__1), .A1 (
          nx35986), .B0 (camera_module_cache_ram_81__1), .B1 (nx36026)) ;
    dffr camera_module_cache_reg_ram_65__1 (.Q (camera_module_cache_ram_65__1), 
         .QB (\$dummy [1074]), .D (nx6183), .CLK (clk), .R (rst)) ;
    mux21_ni ix6184 (.Y (nx6183), .A0 (camera_module_cache_ram_65__1), .A1 (
             nx35144), .S0 (nx35048)) ;
    dffr camera_module_cache_reg_ram_81__1 (.Q (camera_module_cache_ram_81__1), 
         .QB (\$dummy [1075]), .D (nx6173), .CLK (clk), .R (rst)) ;
    mux21_ni ix6174 (.Y (nx6173), .A0 (camera_module_cache_ram_81__1), .A1 (
             nx35146), .S0 (nx35044)) ;
    aoi22 ix28961 (.Y (nx28960), .A0 (camera_module_cache_ram_113__1), .A1 (
          nx36066), .B0 (camera_module_cache_ram_97__1), .B1 (nx36106)) ;
    dffr camera_module_cache_reg_ram_113__1 (.Q (camera_module_cache_ram_113__1)
         , .QB (\$dummy [1076]), .D (nx6153), .CLK (clk), .R (rst)) ;
    mux21_ni ix6154 (.Y (nx6153), .A0 (camera_module_cache_ram_113__1), .A1 (
             nx35146), .S0 (nx35036)) ;
    dffr camera_module_cache_reg_ram_97__1 (.Q (camera_module_cache_ram_97__1), 
         .QB (\$dummy [1077]), .D (nx6163), .CLK (clk), .R (rst)) ;
    mux21_ni ix6164 (.Y (nx6163), .A0 (camera_module_cache_ram_97__1), .A1 (
             nx35146), .S0 (nx35040)) ;
    nand04 ix8469 (.Y (nx8468), .A0 (nx28969), .A1 (nx28977), .A2 (nx28985), .A3 (
           nx28993)) ;
    aoi22 ix28970 (.Y (nx28969), .A0 (camera_module_cache_ram_129__1), .A1 (
          nx36146), .B0 (camera_module_cache_ram_145__1), .B1 (nx36186)) ;
    dffr camera_module_cache_reg_ram_129__1 (.Q (camera_module_cache_ram_129__1)
         , .QB (\$dummy [1078]), .D (nx6143), .CLK (clk), .R (rst)) ;
    mux21_ni ix6144 (.Y (nx6143), .A0 (camera_module_cache_ram_129__1), .A1 (
             nx35146), .S0 (nx35032)) ;
    dffr camera_module_cache_reg_ram_145__1 (.Q (camera_module_cache_ram_145__1)
         , .QB (\$dummy [1079]), .D (nx6133), .CLK (clk), .R (rst)) ;
    mux21_ni ix6134 (.Y (nx6133), .A0 (camera_module_cache_ram_145__1), .A1 (
             nx35146), .S0 (nx35028)) ;
    aoi22 ix28978 (.Y (nx28977), .A0 (camera_module_cache_ram_177__1), .A1 (
          nx36226), .B0 (camera_module_cache_ram_161__1), .B1 (nx36266)) ;
    dffr camera_module_cache_reg_ram_177__1 (.Q (camera_module_cache_ram_177__1)
         , .QB (\$dummy [1080]), .D (nx6113), .CLK (clk), .R (rst)) ;
    mux21_ni ix6114 (.Y (nx6113), .A0 (camera_module_cache_ram_177__1), .A1 (
             nx35146), .S0 (nx35020)) ;
    dffr camera_module_cache_reg_ram_161__1 (.Q (camera_module_cache_ram_161__1)
         , .QB (\$dummy [1081]), .D (nx6123), .CLK (clk), .R (rst)) ;
    mux21_ni ix6124 (.Y (nx6123), .A0 (camera_module_cache_ram_161__1), .A1 (
             nx35146), .S0 (nx35024)) ;
    aoi22 ix28986 (.Y (nx28985), .A0 (camera_module_cache_ram_193__1), .A1 (
          nx36306), .B0 (camera_module_cache_ram_209__1), .B1 (nx36346)) ;
    dffr camera_module_cache_reg_ram_193__1 (.Q (camera_module_cache_ram_193__1)
         , .QB (\$dummy [1082]), .D (nx6103), .CLK (clk), .R (rst)) ;
    mux21_ni ix6104 (.Y (nx6103), .A0 (camera_module_cache_ram_193__1), .A1 (
             nx35148), .S0 (nx35016)) ;
    dffr camera_module_cache_reg_ram_209__1 (.Q (camera_module_cache_ram_209__1)
         , .QB (\$dummy [1083]), .D (nx6093), .CLK (clk), .R (rst)) ;
    mux21_ni ix6094 (.Y (nx6093), .A0 (camera_module_cache_ram_209__1), .A1 (
             nx35148), .S0 (nx35012)) ;
    aoi22 ix28994 (.Y (nx28993), .A0 (camera_module_cache_ram_225__1), .A1 (
          nx36386), .B0 (camera_module_cache_ram_241__1), .B1 (nx36426)) ;
    dffr camera_module_cache_reg_ram_225__1 (.Q (camera_module_cache_ram_225__1)
         , .QB (\$dummy [1084]), .D (nx6083), .CLK (clk), .R (rst)) ;
    mux21_ni ix6084 (.Y (nx6083), .A0 (camera_module_cache_ram_225__1), .A1 (
             nx35148), .S0 (nx35008)) ;
    dffr camera_module_cache_reg_ram_241__1 (.Q (camera_module_cache_ram_241__1)
         , .QB (\$dummy [1085]), .D (nx6073), .CLK (clk), .R (rst)) ;
    mux21_ni ix6074 (.Y (nx6073), .A0 (camera_module_cache_ram_241__1), .A1 (
             nx35148), .S0 (nx35004)) ;
    oai21 ix29002 (.Y (nx29001), .A0 (nx8382), .A1 (nx8304), .B0 (nx36456)) ;
    nand04 ix8383 (.Y (nx8382), .A0 (nx29004), .A1 (nx29012), .A2 (nx29020), .A3 (
           nx29028)) ;
    aoi22 ix29005 (.Y (nx29004), .A0 (camera_module_cache_ram_2__1), .A1 (
          nx35828), .B0 (camera_module_cache_ram_18__1), .B1 (nx35868)) ;
    dffr camera_module_cache_reg_ram_2__1 (.Q (camera_module_cache_ram_2__1), .QB (
         \$dummy [1086]), .D (nx6063), .CLK (clk), .R (rst)) ;
    mux21_ni ix6064 (.Y (nx6063), .A0 (camera_module_cache_ram_2__1), .A1 (
             nx35148), .S0 (nx34994)) ;
    dffr camera_module_cache_reg_ram_18__1 (.Q (camera_module_cache_ram_18__1), 
         .QB (\$dummy [1087]), .D (nx6053), .CLK (clk), .R (rst)) ;
    mux21_ni ix6054 (.Y (nx6053), .A0 (camera_module_cache_ram_18__1), .A1 (
             nx35148), .S0 (nx34990)) ;
    aoi22 ix29013 (.Y (nx29012), .A0 (camera_module_cache_ram_34__1), .A1 (
          nx35908), .B0 (camera_module_cache_ram_50__1), .B1 (nx35948)) ;
    dffr camera_module_cache_reg_ram_34__1 (.Q (camera_module_cache_ram_34__1), 
         .QB (\$dummy [1088]), .D (nx6043), .CLK (clk), .R (rst)) ;
    mux21_ni ix6044 (.Y (nx6043), .A0 (camera_module_cache_ram_34__1), .A1 (
             nx35148), .S0 (nx34986)) ;
    dffr camera_module_cache_reg_ram_50__1 (.Q (camera_module_cache_ram_50__1), 
         .QB (\$dummy [1089]), .D (nx6033), .CLK (clk), .R (rst)) ;
    mux21_ni ix6034 (.Y (nx6033), .A0 (camera_module_cache_ram_50__1), .A1 (
             nx35150), .S0 (nx34982)) ;
    aoi22 ix29021 (.Y (nx29020), .A0 (camera_module_cache_ram_66__1), .A1 (
          nx35988), .B0 (camera_module_cache_ram_82__1), .B1 (nx36028)) ;
    dffr camera_module_cache_reg_ram_66__1 (.Q (camera_module_cache_ram_66__1), 
         .QB (\$dummy [1090]), .D (nx6023), .CLK (clk), .R (rst)) ;
    mux21_ni ix6024 (.Y (nx6023), .A0 (camera_module_cache_ram_66__1), .A1 (
             nx35150), .S0 (nx34978)) ;
    dffr camera_module_cache_reg_ram_82__1 (.Q (camera_module_cache_ram_82__1), 
         .QB (\$dummy [1091]), .D (nx6013), .CLK (clk), .R (rst)) ;
    mux21_ni ix6014 (.Y (nx6013), .A0 (camera_module_cache_ram_82__1), .A1 (
             nx35150), .S0 (nx34974)) ;
    aoi22 ix29029 (.Y (nx29028), .A0 (camera_module_cache_ram_114__1), .A1 (
          nx36068), .B0 (camera_module_cache_ram_98__1), .B1 (nx36108)) ;
    dffr camera_module_cache_reg_ram_114__1 (.Q (camera_module_cache_ram_114__1)
         , .QB (\$dummy [1092]), .D (nx5993), .CLK (clk), .R (rst)) ;
    mux21_ni ix5994 (.Y (nx5993), .A0 (camera_module_cache_ram_114__1), .A1 (
             nx35150), .S0 (nx34966)) ;
    dffr camera_module_cache_reg_ram_98__1 (.Q (camera_module_cache_ram_98__1), 
         .QB (\$dummy [1093]), .D (nx6003), .CLK (clk), .R (rst)) ;
    mux21_ni ix6004 (.Y (nx6003), .A0 (camera_module_cache_ram_98__1), .A1 (
             nx35150), .S0 (nx34970)) ;
    nand04 ix8305 (.Y (nx8304), .A0 (nx29037), .A1 (nx29045), .A2 (nx29053), .A3 (
           nx29061)) ;
    aoi22 ix29038 (.Y (nx29037), .A0 (camera_module_cache_ram_130__1), .A1 (
          nx36148), .B0 (camera_module_cache_ram_146__1), .B1 (nx36188)) ;
    dffr camera_module_cache_reg_ram_130__1 (.Q (camera_module_cache_ram_130__1)
         , .QB (\$dummy [1094]), .D (nx5983), .CLK (clk), .R (rst)) ;
    mux21_ni ix5984 (.Y (nx5983), .A0 (camera_module_cache_ram_130__1), .A1 (
             nx35150), .S0 (nx34962)) ;
    dffr camera_module_cache_reg_ram_146__1 (.Q (camera_module_cache_ram_146__1)
         , .QB (\$dummy [1095]), .D (nx5973), .CLK (clk), .R (rst)) ;
    mux21_ni ix5974 (.Y (nx5973), .A0 (camera_module_cache_ram_146__1), .A1 (
             nx35150), .S0 (nx34958)) ;
    aoi22 ix29046 (.Y (nx29045), .A0 (camera_module_cache_ram_178__1), .A1 (
          nx36228), .B0 (camera_module_cache_ram_162__1), .B1 (nx36268)) ;
    dffr camera_module_cache_reg_ram_178__1 (.Q (camera_module_cache_ram_178__1)
         , .QB (\$dummy [1096]), .D (nx5953), .CLK (clk), .R (rst)) ;
    mux21_ni ix5954 (.Y (nx5953), .A0 (camera_module_cache_ram_178__1), .A1 (
             nx35152), .S0 (nx34950)) ;
    dffr camera_module_cache_reg_ram_162__1 (.Q (camera_module_cache_ram_162__1)
         , .QB (\$dummy [1097]), .D (nx5963), .CLK (clk), .R (rst)) ;
    mux21_ni ix5964 (.Y (nx5963), .A0 (camera_module_cache_ram_162__1), .A1 (
             nx35152), .S0 (nx34954)) ;
    aoi22 ix29054 (.Y (nx29053), .A0 (camera_module_cache_ram_194__1), .A1 (
          nx36308), .B0 (camera_module_cache_ram_210__1), .B1 (nx36348)) ;
    dffr camera_module_cache_reg_ram_194__1 (.Q (camera_module_cache_ram_194__1)
         , .QB (\$dummy [1098]), .D (nx5943), .CLK (clk), .R (rst)) ;
    mux21_ni ix5944 (.Y (nx5943), .A0 (camera_module_cache_ram_194__1), .A1 (
             nx35152), .S0 (nx34946)) ;
    dffr camera_module_cache_reg_ram_210__1 (.Q (camera_module_cache_ram_210__1)
         , .QB (\$dummy [1099]), .D (nx5933), .CLK (clk), .R (rst)) ;
    mux21_ni ix5934 (.Y (nx5933), .A0 (camera_module_cache_ram_210__1), .A1 (
             nx35152), .S0 (nx34942)) ;
    aoi22 ix29062 (.Y (nx29061), .A0 (camera_module_cache_ram_226__1), .A1 (
          nx36388), .B0 (camera_module_cache_ram_242__1), .B1 (nx36428)) ;
    dffr camera_module_cache_reg_ram_226__1 (.Q (camera_module_cache_ram_226__1)
         , .QB (\$dummy [1100]), .D (nx5923), .CLK (clk), .R (rst)) ;
    mux21_ni ix5924 (.Y (nx5923), .A0 (camera_module_cache_ram_226__1), .A1 (
             nx35152), .S0 (nx34938)) ;
    dffr camera_module_cache_reg_ram_242__1 (.Q (camera_module_cache_ram_242__1)
         , .QB (\$dummy [1101]), .D (nx5913), .CLK (clk), .R (rst)) ;
    mux21_ni ix5914 (.Y (nx5913), .A0 (camera_module_cache_ram_242__1), .A1 (
             nx35152), .S0 (nx34934)) ;
    oai21 ix29070 (.Y (nx29069), .A0 (nx8220), .A1 (nx8142), .B0 (nx36460)) ;
    nand04 ix8221 (.Y (nx8220), .A0 (nx29072), .A1 (nx29080), .A2 (nx29088), .A3 (
           nx29096)) ;
    aoi22 ix29073 (.Y (nx29072), .A0 (camera_module_cache_ram_3__1), .A1 (
          nx35828), .B0 (camera_module_cache_ram_19__1), .B1 (nx35868)) ;
    dffr camera_module_cache_reg_ram_3__1 (.Q (camera_module_cache_ram_3__1), .QB (
         \$dummy [1102]), .D (nx5903), .CLK (clk), .R (rst)) ;
    mux21_ni ix5904 (.Y (nx5903), .A0 (camera_module_cache_ram_3__1), .A1 (
             nx35152), .S0 (nx34924)) ;
    dffr camera_module_cache_reg_ram_19__1 (.Q (camera_module_cache_ram_19__1), 
         .QB (\$dummy [1103]), .D (nx5893), .CLK (clk), .R (rst)) ;
    mux21_ni ix5894 (.Y (nx5893), .A0 (camera_module_cache_ram_19__1), .A1 (
             nx35154), .S0 (nx34920)) ;
    aoi22 ix29081 (.Y (nx29080), .A0 (camera_module_cache_ram_35__1), .A1 (
          nx35908), .B0 (camera_module_cache_ram_51__1), .B1 (nx35948)) ;
    dffr camera_module_cache_reg_ram_35__1 (.Q (camera_module_cache_ram_35__1), 
         .QB (\$dummy [1104]), .D (nx5883), .CLK (clk), .R (rst)) ;
    mux21_ni ix5884 (.Y (nx5883), .A0 (camera_module_cache_ram_35__1), .A1 (
             nx35154), .S0 (nx34916)) ;
    dffr camera_module_cache_reg_ram_51__1 (.Q (camera_module_cache_ram_51__1), 
         .QB (\$dummy [1105]), .D (nx5873), .CLK (clk), .R (rst)) ;
    mux21_ni ix5874 (.Y (nx5873), .A0 (camera_module_cache_ram_51__1), .A1 (
             nx35154), .S0 (nx34912)) ;
    aoi22 ix29089 (.Y (nx29088), .A0 (camera_module_cache_ram_67__1), .A1 (
          nx35988), .B0 (camera_module_cache_ram_83__1), .B1 (nx36028)) ;
    dffr camera_module_cache_reg_ram_67__1 (.Q (camera_module_cache_ram_67__1), 
         .QB (\$dummy [1106]), .D (nx5863), .CLK (clk), .R (rst)) ;
    mux21_ni ix5864 (.Y (nx5863), .A0 (camera_module_cache_ram_67__1), .A1 (
             nx35154), .S0 (nx34908)) ;
    dffr camera_module_cache_reg_ram_83__1 (.Q (camera_module_cache_ram_83__1), 
         .QB (\$dummy [1107]), .D (nx5853), .CLK (clk), .R (rst)) ;
    mux21_ni ix5854 (.Y (nx5853), .A0 (camera_module_cache_ram_83__1), .A1 (
             nx35154), .S0 (nx34904)) ;
    aoi22 ix29097 (.Y (nx29096), .A0 (camera_module_cache_ram_115__1), .A1 (
          nx36068), .B0 (camera_module_cache_ram_99__1), .B1 (nx36108)) ;
    dffr camera_module_cache_reg_ram_115__1 (.Q (camera_module_cache_ram_115__1)
         , .QB (\$dummy [1108]), .D (nx5833), .CLK (clk), .R (rst)) ;
    mux21_ni ix5834 (.Y (nx5833), .A0 (camera_module_cache_ram_115__1), .A1 (
             nx35154), .S0 (nx34896)) ;
    dffr camera_module_cache_reg_ram_99__1 (.Q (camera_module_cache_ram_99__1), 
         .QB (\$dummy [1109]), .D (nx5843), .CLK (clk), .R (rst)) ;
    mux21_ni ix5844 (.Y (nx5843), .A0 (camera_module_cache_ram_99__1), .A1 (
             nx35154), .S0 (nx34900)) ;
    nand04 ix8143 (.Y (nx8142), .A0 (nx29105), .A1 (nx29113), .A2 (nx29121), .A3 (
           nx29129)) ;
    aoi22 ix29106 (.Y (nx29105), .A0 (camera_module_cache_ram_131__1), .A1 (
          nx36148), .B0 (camera_module_cache_ram_147__1), .B1 (nx36188)) ;
    dffr camera_module_cache_reg_ram_131__1 (.Q (camera_module_cache_ram_131__1)
         , .QB (\$dummy [1110]), .D (nx5823), .CLK (clk), .R (rst)) ;
    mux21_ni ix5824 (.Y (nx5823), .A0 (camera_module_cache_ram_131__1), .A1 (
             nx35156), .S0 (nx34892)) ;
    dffr camera_module_cache_reg_ram_147__1 (.Q (camera_module_cache_ram_147__1)
         , .QB (\$dummy [1111]), .D (nx5813), .CLK (clk), .R (rst)) ;
    mux21_ni ix5814 (.Y (nx5813), .A0 (camera_module_cache_ram_147__1), .A1 (
             nx35156), .S0 (nx34888)) ;
    aoi22 ix29114 (.Y (nx29113), .A0 (camera_module_cache_ram_179__1), .A1 (
          nx36228), .B0 (camera_module_cache_ram_163__1), .B1 (nx36268)) ;
    dffr camera_module_cache_reg_ram_179__1 (.Q (camera_module_cache_ram_179__1)
         , .QB (\$dummy [1112]), .D (nx5793), .CLK (clk), .R (rst)) ;
    mux21_ni ix5794 (.Y (nx5793), .A0 (camera_module_cache_ram_179__1), .A1 (
             nx35156), .S0 (nx34880)) ;
    dffr camera_module_cache_reg_ram_163__1 (.Q (camera_module_cache_ram_163__1)
         , .QB (\$dummy [1113]), .D (nx5803), .CLK (clk), .R (rst)) ;
    mux21_ni ix5804 (.Y (nx5803), .A0 (camera_module_cache_ram_163__1), .A1 (
             nx35156), .S0 (nx34884)) ;
    aoi22 ix29122 (.Y (nx29121), .A0 (camera_module_cache_ram_195__1), .A1 (
          nx36308), .B0 (camera_module_cache_ram_211__1), .B1 (nx36348)) ;
    dffr camera_module_cache_reg_ram_195__1 (.Q (camera_module_cache_ram_195__1)
         , .QB (\$dummy [1114]), .D (nx5783), .CLK (clk), .R (rst)) ;
    mux21_ni ix5784 (.Y (nx5783), .A0 (camera_module_cache_ram_195__1), .A1 (
             nx35156), .S0 (nx34876)) ;
    dffr camera_module_cache_reg_ram_211__1 (.Q (camera_module_cache_ram_211__1)
         , .QB (\$dummy [1115]), .D (nx5773), .CLK (clk), .R (rst)) ;
    mux21_ni ix5774 (.Y (nx5773), .A0 (camera_module_cache_ram_211__1), .A1 (
             nx35156), .S0 (nx34872)) ;
    aoi22 ix29130 (.Y (nx29129), .A0 (camera_module_cache_ram_227__1), .A1 (
          nx36388), .B0 (camera_module_cache_ram_243__1), .B1 (nx36428)) ;
    dffr camera_module_cache_reg_ram_227__1 (.Q (camera_module_cache_ram_227__1)
         , .QB (\$dummy [1116]), .D (nx5763), .CLK (clk), .R (rst)) ;
    mux21_ni ix5764 (.Y (nx5763), .A0 (camera_module_cache_ram_227__1), .A1 (
             nx35156), .S0 (nx34868)) ;
    dffr camera_module_cache_reg_ram_243__1 (.Q (camera_module_cache_ram_243__1)
         , .QB (\$dummy [1117]), .D (nx5753), .CLK (clk), .R (rst)) ;
    mux21_ni ix5754 (.Y (nx5753), .A0 (camera_module_cache_ram_243__1), .A1 (
             nx35158), .S0 (nx34864)) ;
    nand04 ix8065 (.Y (nx8064), .A0 (nx29138), .A1 (nx29206), .A2 (nx29274), .A3 (
           nx29342)) ;
    oai21 ix29139 (.Y (nx29138), .A0 (nx8054), .A1 (nx7976), .B0 (nx36464)) ;
    nand04 ix8055 (.Y (nx8054), .A0 (nx29141), .A1 (nx29149), .A2 (nx29157), .A3 (
           nx29165)) ;
    aoi22 ix29142 (.Y (nx29141), .A0 (camera_module_cache_ram_4__1), .A1 (
          nx35828), .B0 (camera_module_cache_ram_20__1), .B1 (nx35868)) ;
    dffr camera_module_cache_reg_ram_4__1 (.Q (camera_module_cache_ram_4__1), .QB (
         \$dummy [1118]), .D (nx5743), .CLK (clk), .R (rst)) ;
    mux21_ni ix5744 (.Y (nx5743), .A0 (camera_module_cache_ram_4__1), .A1 (
             nx35158), .S0 (nx34854)) ;
    dffr camera_module_cache_reg_ram_20__1 (.Q (camera_module_cache_ram_20__1), 
         .QB (\$dummy [1119]), .D (nx5733), .CLK (clk), .R (rst)) ;
    mux21_ni ix5734 (.Y (nx5733), .A0 (camera_module_cache_ram_20__1), .A1 (
             nx35158), .S0 (nx34850)) ;
    aoi22 ix29150 (.Y (nx29149), .A0 (camera_module_cache_ram_36__1), .A1 (
          nx35908), .B0 (camera_module_cache_ram_52__1), .B1 (nx35948)) ;
    dffr camera_module_cache_reg_ram_36__1 (.Q (camera_module_cache_ram_36__1), 
         .QB (\$dummy [1120]), .D (nx5723), .CLK (clk), .R (rst)) ;
    mux21_ni ix5724 (.Y (nx5723), .A0 (camera_module_cache_ram_36__1), .A1 (
             nx35158), .S0 (nx34846)) ;
    dffr camera_module_cache_reg_ram_52__1 (.Q (camera_module_cache_ram_52__1), 
         .QB (\$dummy [1121]), .D (nx5713), .CLK (clk), .R (rst)) ;
    mux21_ni ix5714 (.Y (nx5713), .A0 (camera_module_cache_ram_52__1), .A1 (
             nx35158), .S0 (nx34842)) ;
    aoi22 ix29158 (.Y (nx29157), .A0 (camera_module_cache_ram_68__1), .A1 (
          nx35988), .B0 (camera_module_cache_ram_84__1), .B1 (nx36028)) ;
    dffr camera_module_cache_reg_ram_68__1 (.Q (camera_module_cache_ram_68__1), 
         .QB (\$dummy [1122]), .D (nx5703), .CLK (clk), .R (rst)) ;
    mux21_ni ix5704 (.Y (nx5703), .A0 (camera_module_cache_ram_68__1), .A1 (
             nx35158), .S0 (nx34838)) ;
    dffr camera_module_cache_reg_ram_84__1 (.Q (camera_module_cache_ram_84__1), 
         .QB (\$dummy [1123]), .D (nx5693), .CLK (clk), .R (rst)) ;
    mux21_ni ix5694 (.Y (nx5693), .A0 (camera_module_cache_ram_84__1), .A1 (
             nx35158), .S0 (nx34834)) ;
    aoi22 ix29166 (.Y (nx29165), .A0 (camera_module_cache_ram_116__1), .A1 (
          nx36068), .B0 (camera_module_cache_ram_100__1), .B1 (nx36108)) ;
    dffr camera_module_cache_reg_ram_116__1 (.Q (camera_module_cache_ram_116__1)
         , .QB (\$dummy [1124]), .D (nx5673), .CLK (clk), .R (rst)) ;
    mux21_ni ix5674 (.Y (nx5673), .A0 (camera_module_cache_ram_116__1), .A1 (
             nx35160), .S0 (nx34826)) ;
    dffr camera_module_cache_reg_ram_100__1 (.Q (camera_module_cache_ram_100__1)
         , .QB (\$dummy [1125]), .D (nx5683), .CLK (clk), .R (rst)) ;
    mux21_ni ix5684 (.Y (nx5683), .A0 (camera_module_cache_ram_100__1), .A1 (
             nx35160), .S0 (nx34830)) ;
    nand04 ix7977 (.Y (nx7976), .A0 (nx29174), .A1 (nx29182), .A2 (nx29190), .A3 (
           nx29198)) ;
    aoi22 ix29175 (.Y (nx29174), .A0 (camera_module_cache_ram_132__1), .A1 (
          nx36148), .B0 (camera_module_cache_ram_148__1), .B1 (nx36188)) ;
    dffr camera_module_cache_reg_ram_132__1 (.Q (camera_module_cache_ram_132__1)
         , .QB (\$dummy [1126]), .D (nx5663), .CLK (clk), .R (rst)) ;
    mux21_ni ix5664 (.Y (nx5663), .A0 (camera_module_cache_ram_132__1), .A1 (
             nx35160), .S0 (nx34822)) ;
    dffr camera_module_cache_reg_ram_148__1 (.Q (camera_module_cache_ram_148__1)
         , .QB (\$dummy [1127]), .D (nx5653), .CLK (clk), .R (rst)) ;
    mux21_ni ix5654 (.Y (nx5653), .A0 (camera_module_cache_ram_148__1), .A1 (
             nx35160), .S0 (nx34818)) ;
    aoi22 ix29183 (.Y (nx29182), .A0 (camera_module_cache_ram_180__1), .A1 (
          nx36228), .B0 (camera_module_cache_ram_164__1), .B1 (nx36268)) ;
    dffr camera_module_cache_reg_ram_180__1 (.Q (camera_module_cache_ram_180__1)
         , .QB (\$dummy [1128]), .D (nx5633), .CLK (clk), .R (rst)) ;
    mux21_ni ix5634 (.Y (nx5633), .A0 (camera_module_cache_ram_180__1), .A1 (
             nx35160), .S0 (nx34810)) ;
    dffr camera_module_cache_reg_ram_164__1 (.Q (camera_module_cache_ram_164__1)
         , .QB (\$dummy [1129]), .D (nx5643), .CLK (clk), .R (rst)) ;
    mux21_ni ix5644 (.Y (nx5643), .A0 (camera_module_cache_ram_164__1), .A1 (
             nx35160), .S0 (nx34814)) ;
    aoi22 ix29191 (.Y (nx29190), .A0 (camera_module_cache_ram_196__1), .A1 (
          nx36308), .B0 (camera_module_cache_ram_212__1), .B1 (nx36348)) ;
    dffr camera_module_cache_reg_ram_196__1 (.Q (camera_module_cache_ram_196__1)
         , .QB (\$dummy [1130]), .D (nx5623), .CLK (clk), .R (rst)) ;
    mux21_ni ix5624 (.Y (nx5623), .A0 (camera_module_cache_ram_196__1), .A1 (
             nx35160), .S0 (nx34806)) ;
    dffr camera_module_cache_reg_ram_212__1 (.Q (camera_module_cache_ram_212__1)
         , .QB (\$dummy [1131]), .D (nx5613), .CLK (clk), .R (rst)) ;
    mux21_ni ix5614 (.Y (nx5613), .A0 (camera_module_cache_ram_212__1), .A1 (
             nx35162), .S0 (nx34802)) ;
    aoi22 ix29199 (.Y (nx29198), .A0 (camera_module_cache_ram_228__1), .A1 (
          nx36388), .B0 (camera_module_cache_ram_244__1), .B1 (nx36428)) ;
    dffr camera_module_cache_reg_ram_228__1 (.Q (camera_module_cache_ram_228__1)
         , .QB (\$dummy [1132]), .D (nx5603), .CLK (clk), .R (rst)) ;
    mux21_ni ix5604 (.Y (nx5603), .A0 (camera_module_cache_ram_228__1), .A1 (
             nx35162), .S0 (nx34798)) ;
    dffr camera_module_cache_reg_ram_244__1 (.Q (camera_module_cache_ram_244__1)
         , .QB (\$dummy [1133]), .D (nx5593), .CLK (clk), .R (rst)) ;
    mux21_ni ix5594 (.Y (nx5593), .A0 (camera_module_cache_ram_244__1), .A1 (
             nx35162), .S0 (nx34794)) ;
    oai21 ix29207 (.Y (nx29206), .A0 (nx7892), .A1 (nx7814), .B0 (nx36468)) ;
    nand04 ix7893 (.Y (nx7892), .A0 (nx29209), .A1 (nx29217), .A2 (nx29225), .A3 (
           nx29233)) ;
    aoi22 ix29210 (.Y (nx29209), .A0 (camera_module_cache_ram_5__1), .A1 (
          nx35828), .B0 (camera_module_cache_ram_21__1), .B1 (nx35868)) ;
    dffr camera_module_cache_reg_ram_5__1 (.Q (camera_module_cache_ram_5__1), .QB (
         \$dummy [1134]), .D (nx5583), .CLK (clk), .R (rst)) ;
    mux21_ni ix5584 (.Y (nx5583), .A0 (camera_module_cache_ram_5__1), .A1 (
             nx35162), .S0 (nx34784)) ;
    dffr camera_module_cache_reg_ram_21__1 (.Q (camera_module_cache_ram_21__1), 
         .QB (\$dummy [1135]), .D (nx5573), .CLK (clk), .R (rst)) ;
    mux21_ni ix5574 (.Y (nx5573), .A0 (camera_module_cache_ram_21__1), .A1 (
             nx35162), .S0 (nx34780)) ;
    aoi22 ix29218 (.Y (nx29217), .A0 (camera_module_cache_ram_37__1), .A1 (
          nx35908), .B0 (camera_module_cache_ram_53__1), .B1 (nx35948)) ;
    dffr camera_module_cache_reg_ram_37__1 (.Q (camera_module_cache_ram_37__1), 
         .QB (\$dummy [1136]), .D (nx5563), .CLK (clk), .R (rst)) ;
    mux21_ni ix5564 (.Y (nx5563), .A0 (camera_module_cache_ram_37__1), .A1 (
             nx35162), .S0 (nx34776)) ;
    dffr camera_module_cache_reg_ram_53__1 (.Q (camera_module_cache_ram_53__1), 
         .QB (\$dummy [1137]), .D (nx5553), .CLK (clk), .R (rst)) ;
    mux21_ni ix5554 (.Y (nx5553), .A0 (camera_module_cache_ram_53__1), .A1 (
             nx35162), .S0 (nx34772)) ;
    aoi22 ix29226 (.Y (nx29225), .A0 (camera_module_cache_ram_69__1), .A1 (
          nx35988), .B0 (camera_module_cache_ram_85__1), .B1 (nx36028)) ;
    dffr camera_module_cache_reg_ram_69__1 (.Q (camera_module_cache_ram_69__1), 
         .QB (\$dummy [1138]), .D (nx5543), .CLK (clk), .R (rst)) ;
    mux21_ni ix5544 (.Y (nx5543), .A0 (camera_module_cache_ram_69__1), .A1 (
             nx35164), .S0 (nx34768)) ;
    dffr camera_module_cache_reg_ram_85__1 (.Q (camera_module_cache_ram_85__1), 
         .QB (\$dummy [1139]), .D (nx5533), .CLK (clk), .R (rst)) ;
    mux21_ni ix5534 (.Y (nx5533), .A0 (camera_module_cache_ram_85__1), .A1 (
             nx35164), .S0 (nx34764)) ;
    aoi22 ix29234 (.Y (nx29233), .A0 (camera_module_cache_ram_117__1), .A1 (
          nx36068), .B0 (camera_module_cache_ram_101__1), .B1 (nx36108)) ;
    dffr camera_module_cache_reg_ram_117__1 (.Q (camera_module_cache_ram_117__1)
         , .QB (\$dummy [1140]), .D (nx5513), .CLK (clk), .R (rst)) ;
    mux21_ni ix5514 (.Y (nx5513), .A0 (camera_module_cache_ram_117__1), .A1 (
             nx35164), .S0 (nx34756)) ;
    dffr camera_module_cache_reg_ram_101__1 (.Q (camera_module_cache_ram_101__1)
         , .QB (\$dummy [1141]), .D (nx5523), .CLK (clk), .R (rst)) ;
    mux21_ni ix5524 (.Y (nx5523), .A0 (camera_module_cache_ram_101__1), .A1 (
             nx35164), .S0 (nx34760)) ;
    nand04 ix7815 (.Y (nx7814), .A0 (nx29242), .A1 (nx29250), .A2 (nx29258), .A3 (
           nx29266)) ;
    aoi22 ix29243 (.Y (nx29242), .A0 (camera_module_cache_ram_133__1), .A1 (
          nx36148), .B0 (camera_module_cache_ram_149__1), .B1 (nx36188)) ;
    dffr camera_module_cache_reg_ram_133__1 (.Q (camera_module_cache_ram_133__1)
         , .QB (\$dummy [1142]), .D (nx5503), .CLK (clk), .R (rst)) ;
    mux21_ni ix5504 (.Y (nx5503), .A0 (camera_module_cache_ram_133__1), .A1 (
             nx35164), .S0 (nx34752)) ;
    dffr camera_module_cache_reg_ram_149__1 (.Q (camera_module_cache_ram_149__1)
         , .QB (\$dummy [1143]), .D (nx5493), .CLK (clk), .R (rst)) ;
    mux21_ni ix5494 (.Y (nx5493), .A0 (camera_module_cache_ram_149__1), .A1 (
             nx35164), .S0 (nx34748)) ;
    aoi22 ix29251 (.Y (nx29250), .A0 (camera_module_cache_ram_181__1), .A1 (
          nx36228), .B0 (camera_module_cache_ram_165__1), .B1 (nx36268)) ;
    dffr camera_module_cache_reg_ram_181__1 (.Q (camera_module_cache_ram_181__1)
         , .QB (\$dummy [1144]), .D (nx5473), .CLK (clk), .R (rst)) ;
    mux21_ni ix5474 (.Y (nx5473), .A0 (camera_module_cache_ram_181__1), .A1 (
             nx35164), .S0 (nx34740)) ;
    dffr camera_module_cache_reg_ram_165__1 (.Q (camera_module_cache_ram_165__1)
         , .QB (\$dummy [1145]), .D (nx5483), .CLK (clk), .R (rst)) ;
    mux21_ni ix5484 (.Y (nx5483), .A0 (camera_module_cache_ram_165__1), .A1 (
             nx35166), .S0 (nx34744)) ;
    aoi22 ix29259 (.Y (nx29258), .A0 (camera_module_cache_ram_197__1), .A1 (
          nx36308), .B0 (camera_module_cache_ram_213__1), .B1 (nx36348)) ;
    dffr camera_module_cache_reg_ram_197__1 (.Q (camera_module_cache_ram_197__1)
         , .QB (\$dummy [1146]), .D (nx5463), .CLK (clk), .R (rst)) ;
    mux21_ni ix5464 (.Y (nx5463), .A0 (camera_module_cache_ram_197__1), .A1 (
             nx35166), .S0 (nx34736)) ;
    dffr camera_module_cache_reg_ram_213__1 (.Q (camera_module_cache_ram_213__1)
         , .QB (\$dummy [1147]), .D (nx5453), .CLK (clk), .R (rst)) ;
    mux21_ni ix5454 (.Y (nx5453), .A0 (camera_module_cache_ram_213__1), .A1 (
             nx35166), .S0 (nx34732)) ;
    aoi22 ix29267 (.Y (nx29266), .A0 (camera_module_cache_ram_229__1), .A1 (
          nx36388), .B0 (camera_module_cache_ram_245__1), .B1 (nx36428)) ;
    dffr camera_module_cache_reg_ram_229__1 (.Q (camera_module_cache_ram_229__1)
         , .QB (\$dummy [1148]), .D (nx5443), .CLK (clk), .R (rst)) ;
    mux21_ni ix5444 (.Y (nx5443), .A0 (camera_module_cache_ram_229__1), .A1 (
             nx35166), .S0 (nx34728)) ;
    dffr camera_module_cache_reg_ram_245__1 (.Q (camera_module_cache_ram_245__1)
         , .QB (\$dummy [1149]), .D (nx5433), .CLK (clk), .R (rst)) ;
    mux21_ni ix5434 (.Y (nx5433), .A0 (camera_module_cache_ram_245__1), .A1 (
             nx35166), .S0 (nx34724)) ;
    oai21 ix29275 (.Y (nx29274), .A0 (nx7728), .A1 (nx7650), .B0 (nx36472)) ;
    nand04 ix7729 (.Y (nx7728), .A0 (nx29277), .A1 (nx29285), .A2 (nx29293), .A3 (
           nx29301)) ;
    aoi22 ix29278 (.Y (nx29277), .A0 (camera_module_cache_ram_6__1), .A1 (
          nx35828), .B0 (camera_module_cache_ram_22__1), .B1 (nx35868)) ;
    dffr camera_module_cache_reg_ram_6__1 (.Q (camera_module_cache_ram_6__1), .QB (
         \$dummy [1150]), .D (nx5423), .CLK (clk), .R (rst)) ;
    mux21_ni ix5424 (.Y (nx5423), .A0 (camera_module_cache_ram_6__1), .A1 (
             nx35166), .S0 (nx34714)) ;
    dffr camera_module_cache_reg_ram_22__1 (.Q (camera_module_cache_ram_22__1), 
         .QB (\$dummy [1151]), .D (nx5413), .CLK (clk), .R (rst)) ;
    mux21_ni ix5414 (.Y (nx5413), .A0 (camera_module_cache_ram_22__1), .A1 (
             nx35166), .S0 (nx34710)) ;
    aoi22 ix29286 (.Y (nx29285), .A0 (camera_module_cache_ram_38__1), .A1 (
          nx35908), .B0 (camera_module_cache_ram_54__1), .B1 (nx35948)) ;
    dffr camera_module_cache_reg_ram_38__1 (.Q (camera_module_cache_ram_38__1), 
         .QB (\$dummy [1152]), .D (nx5403), .CLK (clk), .R (rst)) ;
    mux21_ni ix5404 (.Y (nx5403), .A0 (camera_module_cache_ram_38__1), .A1 (
             nx35168), .S0 (nx34706)) ;
    dffr camera_module_cache_reg_ram_54__1 (.Q (camera_module_cache_ram_54__1), 
         .QB (\$dummy [1153]), .D (nx5393), .CLK (clk), .R (rst)) ;
    mux21_ni ix5394 (.Y (nx5393), .A0 (camera_module_cache_ram_54__1), .A1 (
             nx35168), .S0 (nx34702)) ;
    aoi22 ix29294 (.Y (nx29293), .A0 (camera_module_cache_ram_70__1), .A1 (
          nx35988), .B0 (camera_module_cache_ram_86__1), .B1 (nx36028)) ;
    dffr camera_module_cache_reg_ram_70__1 (.Q (camera_module_cache_ram_70__1), 
         .QB (\$dummy [1154]), .D (nx5383), .CLK (clk), .R (rst)) ;
    mux21_ni ix5384 (.Y (nx5383), .A0 (camera_module_cache_ram_70__1), .A1 (
             nx35168), .S0 (nx34698)) ;
    dffr camera_module_cache_reg_ram_86__1 (.Q (camera_module_cache_ram_86__1), 
         .QB (\$dummy [1155]), .D (nx5373), .CLK (clk), .R (rst)) ;
    mux21_ni ix5374 (.Y (nx5373), .A0 (camera_module_cache_ram_86__1), .A1 (
             nx35168), .S0 (nx34694)) ;
    aoi22 ix29302 (.Y (nx29301), .A0 (camera_module_cache_ram_118__1), .A1 (
          nx36068), .B0 (camera_module_cache_ram_102__1), .B1 (nx36108)) ;
    dffr camera_module_cache_reg_ram_118__1 (.Q (camera_module_cache_ram_118__1)
         , .QB (\$dummy [1156]), .D (nx5353), .CLK (clk), .R (rst)) ;
    mux21_ni ix5354 (.Y (nx5353), .A0 (camera_module_cache_ram_118__1), .A1 (
             nx35168), .S0 (nx34686)) ;
    dffr camera_module_cache_reg_ram_102__1 (.Q (camera_module_cache_ram_102__1)
         , .QB (\$dummy [1157]), .D (nx5363), .CLK (clk), .R (rst)) ;
    mux21_ni ix5364 (.Y (nx5363), .A0 (camera_module_cache_ram_102__1), .A1 (
             nx35168), .S0 (nx34690)) ;
    nand04 ix7651 (.Y (nx7650), .A0 (nx29310), .A1 (nx29318), .A2 (nx29326), .A3 (
           nx29334)) ;
    aoi22 ix29311 (.Y (nx29310), .A0 (camera_module_cache_ram_134__1), .A1 (
          nx36148), .B0 (camera_module_cache_ram_150__1), .B1 (nx36188)) ;
    dffr camera_module_cache_reg_ram_134__1 (.Q (camera_module_cache_ram_134__1)
         , .QB (\$dummy [1158]), .D (nx5343), .CLK (clk), .R (rst)) ;
    mux21_ni ix5344 (.Y (nx5343), .A0 (camera_module_cache_ram_134__1), .A1 (
             nx35168), .S0 (nx34682)) ;
    dffr camera_module_cache_reg_ram_150__1 (.Q (camera_module_cache_ram_150__1)
         , .QB (\$dummy [1159]), .D (nx5333), .CLK (clk), .R (rst)) ;
    mux21_ni ix5334 (.Y (nx5333), .A0 (camera_module_cache_ram_150__1), .A1 (
             nx35170), .S0 (nx34678)) ;
    aoi22 ix29319 (.Y (nx29318), .A0 (camera_module_cache_ram_182__1), .A1 (
          nx36228), .B0 (camera_module_cache_ram_166__1), .B1 (nx36268)) ;
    dffr camera_module_cache_reg_ram_182__1 (.Q (camera_module_cache_ram_182__1)
         , .QB (\$dummy [1160]), .D (nx5313), .CLK (clk), .R (rst)) ;
    mux21_ni ix5314 (.Y (nx5313), .A0 (camera_module_cache_ram_182__1), .A1 (
             nx35170), .S0 (nx34670)) ;
    dffr camera_module_cache_reg_ram_166__1 (.Q (camera_module_cache_ram_166__1)
         , .QB (\$dummy [1161]), .D (nx5323), .CLK (clk), .R (rst)) ;
    mux21_ni ix5324 (.Y (nx5323), .A0 (camera_module_cache_ram_166__1), .A1 (
             nx35170), .S0 (nx34674)) ;
    aoi22 ix29327 (.Y (nx29326), .A0 (camera_module_cache_ram_198__1), .A1 (
          nx36308), .B0 (camera_module_cache_ram_214__1), .B1 (nx36348)) ;
    dffr camera_module_cache_reg_ram_198__1 (.Q (camera_module_cache_ram_198__1)
         , .QB (\$dummy [1162]), .D (nx5303), .CLK (clk), .R (rst)) ;
    mux21_ni ix5304 (.Y (nx5303), .A0 (camera_module_cache_ram_198__1), .A1 (
             nx35170), .S0 (nx34666)) ;
    dffr camera_module_cache_reg_ram_214__1 (.Q (camera_module_cache_ram_214__1)
         , .QB (\$dummy [1163]), .D (nx5293), .CLK (clk), .R (rst)) ;
    mux21_ni ix5294 (.Y (nx5293), .A0 (camera_module_cache_ram_214__1), .A1 (
             nx35170), .S0 (nx34662)) ;
    aoi22 ix29335 (.Y (nx29334), .A0 (camera_module_cache_ram_230__1), .A1 (
          nx36388), .B0 (camera_module_cache_ram_246__1), .B1 (nx36428)) ;
    dffr camera_module_cache_reg_ram_230__1 (.Q (camera_module_cache_ram_230__1)
         , .QB (\$dummy [1164]), .D (nx5283), .CLK (clk), .R (rst)) ;
    mux21_ni ix5284 (.Y (nx5283), .A0 (camera_module_cache_ram_230__1), .A1 (
             nx35170), .S0 (nx34658)) ;
    dffr camera_module_cache_reg_ram_246__1 (.Q (camera_module_cache_ram_246__1)
         , .QB (\$dummy [1165]), .D (nx5273), .CLK (clk), .R (rst)) ;
    mux21_ni ix5274 (.Y (nx5273), .A0 (camera_module_cache_ram_246__1), .A1 (
             nx35170), .S0 (nx34654)) ;
    oai21 ix29343 (.Y (nx29342), .A0 (nx7566), .A1 (nx7488), .B0 (nx36476)) ;
    nand04 ix7567 (.Y (nx7566), .A0 (nx29345), .A1 (nx29353), .A2 (nx29361), .A3 (
           nx29369)) ;
    aoi22 ix29346 (.Y (nx29345), .A0 (camera_module_cache_ram_7__1), .A1 (
          nx35828), .B0 (camera_module_cache_ram_23__1), .B1 (nx35868)) ;
    dffr camera_module_cache_reg_ram_7__1 (.Q (camera_module_cache_ram_7__1), .QB (
         \$dummy [1166]), .D (nx5263), .CLK (clk), .R (rst)) ;
    mux21_ni ix5264 (.Y (nx5263), .A0 (camera_module_cache_ram_7__1), .A1 (
             nx35172), .S0 (nx34644)) ;
    dffr camera_module_cache_reg_ram_23__1 (.Q (camera_module_cache_ram_23__1), 
         .QB (\$dummy [1167]), .D (nx5253), .CLK (clk), .R (rst)) ;
    mux21_ni ix5254 (.Y (nx5253), .A0 (camera_module_cache_ram_23__1), .A1 (
             nx35172), .S0 (nx34640)) ;
    aoi22 ix29354 (.Y (nx29353), .A0 (camera_module_cache_ram_39__1), .A1 (
          nx35908), .B0 (camera_module_cache_ram_55__1), .B1 (nx35948)) ;
    dffr camera_module_cache_reg_ram_39__1 (.Q (camera_module_cache_ram_39__1), 
         .QB (\$dummy [1168]), .D (nx5243), .CLK (clk), .R (rst)) ;
    mux21_ni ix5244 (.Y (nx5243), .A0 (camera_module_cache_ram_39__1), .A1 (
             nx35172), .S0 (nx34636)) ;
    dffr camera_module_cache_reg_ram_55__1 (.Q (camera_module_cache_ram_55__1), 
         .QB (\$dummy [1169]), .D (nx5233), .CLK (clk), .R (rst)) ;
    mux21_ni ix5234 (.Y (nx5233), .A0 (camera_module_cache_ram_55__1), .A1 (
             nx35172), .S0 (nx34632)) ;
    aoi22 ix29362 (.Y (nx29361), .A0 (camera_module_cache_ram_71__1), .A1 (
          nx35988), .B0 (camera_module_cache_ram_87__1), .B1 (nx36028)) ;
    dffr camera_module_cache_reg_ram_71__1 (.Q (camera_module_cache_ram_71__1), 
         .QB (\$dummy [1170]), .D (nx5223), .CLK (clk), .R (rst)) ;
    mux21_ni ix5224 (.Y (nx5223), .A0 (camera_module_cache_ram_71__1), .A1 (
             nx35172), .S0 (nx34628)) ;
    dffr camera_module_cache_reg_ram_87__1 (.Q (camera_module_cache_ram_87__1), 
         .QB (\$dummy [1171]), .D (nx5213), .CLK (clk), .R (rst)) ;
    mux21_ni ix5214 (.Y (nx5213), .A0 (camera_module_cache_ram_87__1), .A1 (
             nx35172), .S0 (nx34624)) ;
    aoi22 ix29370 (.Y (nx29369), .A0 (camera_module_cache_ram_119__1), .A1 (
          nx36068), .B0 (camera_module_cache_ram_103__1), .B1 (nx36108)) ;
    dffr camera_module_cache_reg_ram_119__1 (.Q (camera_module_cache_ram_119__1)
         , .QB (\$dummy [1172]), .D (nx5193), .CLK (clk), .R (rst)) ;
    mux21_ni ix5194 (.Y (nx5193), .A0 (camera_module_cache_ram_119__1), .A1 (
             nx35172), .S0 (nx34616)) ;
    dffr camera_module_cache_reg_ram_103__1 (.Q (camera_module_cache_ram_103__1)
         , .QB (\$dummy [1173]), .D (nx5203), .CLK (clk), .R (rst)) ;
    mux21_ni ix5204 (.Y (nx5203), .A0 (camera_module_cache_ram_103__1), .A1 (
             nx35174), .S0 (nx34620)) ;
    nand04 ix7489 (.Y (nx7488), .A0 (nx29378), .A1 (nx29386), .A2 (nx29394), .A3 (
           nx29402)) ;
    aoi22 ix29379 (.Y (nx29378), .A0 (camera_module_cache_ram_135__1), .A1 (
          nx36148), .B0 (camera_module_cache_ram_151__1), .B1 (nx36188)) ;
    dffr camera_module_cache_reg_ram_135__1 (.Q (camera_module_cache_ram_135__1)
         , .QB (\$dummy [1174]), .D (nx5183), .CLK (clk), .R (rst)) ;
    mux21_ni ix5184 (.Y (nx5183), .A0 (camera_module_cache_ram_135__1), .A1 (
             nx35174), .S0 (nx34612)) ;
    dffr camera_module_cache_reg_ram_151__1 (.Q (camera_module_cache_ram_151__1)
         , .QB (\$dummy [1175]), .D (nx5173), .CLK (clk), .R (rst)) ;
    mux21_ni ix5174 (.Y (nx5173), .A0 (camera_module_cache_ram_151__1), .A1 (
             nx35174), .S0 (nx34608)) ;
    aoi22 ix29387 (.Y (nx29386), .A0 (camera_module_cache_ram_183__1), .A1 (
          nx36228), .B0 (camera_module_cache_ram_167__1), .B1 (nx36268)) ;
    dffr camera_module_cache_reg_ram_183__1 (.Q (camera_module_cache_ram_183__1)
         , .QB (\$dummy [1176]), .D (nx5153), .CLK (clk), .R (rst)) ;
    mux21_ni ix5154 (.Y (nx5153), .A0 (camera_module_cache_ram_183__1), .A1 (
             nx35174), .S0 (nx34600)) ;
    dffr camera_module_cache_reg_ram_167__1 (.Q (camera_module_cache_ram_167__1)
         , .QB (\$dummy [1177]), .D (nx5163), .CLK (clk), .R (rst)) ;
    mux21_ni ix5164 (.Y (nx5163), .A0 (camera_module_cache_ram_167__1), .A1 (
             nx35174), .S0 (nx34604)) ;
    aoi22 ix29395 (.Y (nx29394), .A0 (camera_module_cache_ram_199__1), .A1 (
          nx36308), .B0 (camera_module_cache_ram_215__1), .B1 (nx36348)) ;
    dffr camera_module_cache_reg_ram_199__1 (.Q (camera_module_cache_ram_199__1)
         , .QB (\$dummy [1178]), .D (nx5143), .CLK (clk), .R (rst)) ;
    mux21_ni ix5144 (.Y (nx5143), .A0 (camera_module_cache_ram_199__1), .A1 (
             nx35174), .S0 (nx34596)) ;
    dffr camera_module_cache_reg_ram_215__1 (.Q (camera_module_cache_ram_215__1)
         , .QB (\$dummy [1179]), .D (nx5133), .CLK (clk), .R (rst)) ;
    mux21_ni ix5134 (.Y (nx5133), .A0 (camera_module_cache_ram_215__1), .A1 (
             nx35174), .S0 (nx34592)) ;
    aoi22 ix29403 (.Y (nx29402), .A0 (camera_module_cache_ram_231__1), .A1 (
          nx36388), .B0 (camera_module_cache_ram_247__1), .B1 (nx36428)) ;
    dffr camera_module_cache_reg_ram_231__1 (.Q (camera_module_cache_ram_231__1)
         , .QB (\$dummy [1180]), .D (nx5123), .CLK (clk), .R (rst)) ;
    mux21_ni ix5124 (.Y (nx5123), .A0 (camera_module_cache_ram_231__1), .A1 (
             nx35176), .S0 (nx34588)) ;
    dffr camera_module_cache_reg_ram_247__1 (.Q (camera_module_cache_ram_247__1)
         , .QB (\$dummy [1181]), .D (nx5113), .CLK (clk), .R (rst)) ;
    mux21_ni ix5114 (.Y (nx5113), .A0 (camera_module_cache_ram_247__1), .A1 (
             nx35176), .S0 (nx34584)) ;
    nand04 ix7409 (.Y (nx7408), .A0 (nx29411), .A1 (nx29479), .A2 (nx29547), .A3 (
           nx29615)) ;
    oai21 ix29412 (.Y (nx29411), .A0 (nx7398), .A1 (nx7320), .B0 (nx36480)) ;
    nand04 ix7399 (.Y (nx7398), .A0 (nx29414), .A1 (nx29422), .A2 (nx29430), .A3 (
           nx29438)) ;
    aoi22 ix29415 (.Y (nx29414), .A0 (camera_module_cache_ram_8__1), .A1 (
          nx35828), .B0 (camera_module_cache_ram_24__1), .B1 (nx35868)) ;
    dffr camera_module_cache_reg_ram_8__1 (.Q (camera_module_cache_ram_8__1), .QB (
         \$dummy [1182]), .D (nx5103), .CLK (clk), .R (rst)) ;
    mux21_ni ix5104 (.Y (nx5103), .A0 (camera_module_cache_ram_8__1), .A1 (
             nx35176), .S0 (nx34574)) ;
    dffr camera_module_cache_reg_ram_24__1 (.Q (camera_module_cache_ram_24__1), 
         .QB (\$dummy [1183]), .D (nx5093), .CLK (clk), .R (rst)) ;
    mux21_ni ix5094 (.Y (nx5093), .A0 (camera_module_cache_ram_24__1), .A1 (
             nx35176), .S0 (nx34570)) ;
    aoi22 ix29423 (.Y (nx29422), .A0 (camera_module_cache_ram_40__1), .A1 (
          nx35908), .B0 (camera_module_cache_ram_56__1), .B1 (nx35948)) ;
    dffr camera_module_cache_reg_ram_40__1 (.Q (camera_module_cache_ram_40__1), 
         .QB (\$dummy [1184]), .D (nx5083), .CLK (clk), .R (rst)) ;
    mux21_ni ix5084 (.Y (nx5083), .A0 (camera_module_cache_ram_40__1), .A1 (
             nx35176), .S0 (nx34566)) ;
    dffr camera_module_cache_reg_ram_56__1 (.Q (camera_module_cache_ram_56__1), 
         .QB (\$dummy [1185]), .D (nx5073), .CLK (clk), .R (rst)) ;
    mux21_ni ix5074 (.Y (nx5073), .A0 (camera_module_cache_ram_56__1), .A1 (
             nx35176), .S0 (nx34562)) ;
    aoi22 ix29431 (.Y (nx29430), .A0 (camera_module_cache_ram_72__1), .A1 (
          nx35988), .B0 (camera_module_cache_ram_88__1), .B1 (nx36028)) ;
    dffr camera_module_cache_reg_ram_72__1 (.Q (camera_module_cache_ram_72__1), 
         .QB (\$dummy [1186]), .D (nx5063), .CLK (clk), .R (rst)) ;
    mux21_ni ix5064 (.Y (nx5063), .A0 (camera_module_cache_ram_72__1), .A1 (
             nx35176), .S0 (nx34558)) ;
    dffr camera_module_cache_reg_ram_88__1 (.Q (camera_module_cache_ram_88__1), 
         .QB (\$dummy [1187]), .D (nx5053), .CLK (clk), .R (rst)) ;
    mux21_ni ix5054 (.Y (nx5053), .A0 (camera_module_cache_ram_88__1), .A1 (
             nx35178), .S0 (nx34554)) ;
    aoi22 ix29439 (.Y (nx29438), .A0 (camera_module_cache_ram_120__1), .A1 (
          nx36068), .B0 (camera_module_cache_ram_104__1), .B1 (nx36108)) ;
    dffr camera_module_cache_reg_ram_120__1 (.Q (camera_module_cache_ram_120__1)
         , .QB (\$dummy [1188]), .D (nx5033), .CLK (clk), .R (rst)) ;
    mux21_ni ix5034 (.Y (nx5033), .A0 (camera_module_cache_ram_120__1), .A1 (
             nx35178), .S0 (nx34546)) ;
    dffr camera_module_cache_reg_ram_104__1 (.Q (camera_module_cache_ram_104__1)
         , .QB (\$dummy [1189]), .D (nx5043), .CLK (clk), .R (rst)) ;
    mux21_ni ix5044 (.Y (nx5043), .A0 (camera_module_cache_ram_104__1), .A1 (
             nx35178), .S0 (nx34550)) ;
    nand04 ix7321 (.Y (nx7320), .A0 (nx29447), .A1 (nx29455), .A2 (nx29463), .A3 (
           nx29471)) ;
    aoi22 ix29448 (.Y (nx29447), .A0 (camera_module_cache_ram_136__1), .A1 (
          nx36148), .B0 (camera_module_cache_ram_152__1), .B1 (nx36188)) ;
    dffr camera_module_cache_reg_ram_136__1 (.Q (camera_module_cache_ram_136__1)
         , .QB (\$dummy [1190]), .D (nx5023), .CLK (clk), .R (rst)) ;
    mux21_ni ix5024 (.Y (nx5023), .A0 (camera_module_cache_ram_136__1), .A1 (
             nx35178), .S0 (nx34542)) ;
    dffr camera_module_cache_reg_ram_152__1 (.Q (camera_module_cache_ram_152__1)
         , .QB (\$dummy [1191]), .D (nx5013), .CLK (clk), .R (rst)) ;
    mux21_ni ix5014 (.Y (nx5013), .A0 (camera_module_cache_ram_152__1), .A1 (
             nx35178), .S0 (nx34538)) ;
    aoi22 ix29456 (.Y (nx29455), .A0 (camera_module_cache_ram_184__1), .A1 (
          nx36228), .B0 (camera_module_cache_ram_168__1), .B1 (nx36268)) ;
    dffr camera_module_cache_reg_ram_184__1 (.Q (camera_module_cache_ram_184__1)
         , .QB (\$dummy [1192]), .D (nx4993), .CLK (clk), .R (rst)) ;
    mux21_ni ix4994 (.Y (nx4993), .A0 (camera_module_cache_ram_184__1), .A1 (
             nx35178), .S0 (nx34530)) ;
    dffr camera_module_cache_reg_ram_168__1 (.Q (camera_module_cache_ram_168__1)
         , .QB (\$dummy [1193]), .D (nx5003), .CLK (clk), .R (rst)) ;
    mux21_ni ix5004 (.Y (nx5003), .A0 (camera_module_cache_ram_168__1), .A1 (
             nx35178), .S0 (nx34534)) ;
    aoi22 ix29464 (.Y (nx29463), .A0 (camera_module_cache_ram_200__1), .A1 (
          nx36308), .B0 (camera_module_cache_ram_216__1), .B1 (nx36348)) ;
    dffr camera_module_cache_reg_ram_200__1 (.Q (camera_module_cache_ram_200__1)
         , .QB (\$dummy [1194]), .D (nx4983), .CLK (clk), .R (rst)) ;
    mux21_ni ix4984 (.Y (nx4983), .A0 (camera_module_cache_ram_200__1), .A1 (
             nx35180), .S0 (nx34526)) ;
    dffr camera_module_cache_reg_ram_216__1 (.Q (camera_module_cache_ram_216__1)
         , .QB (\$dummy [1195]), .D (nx4973), .CLK (clk), .R (rst)) ;
    mux21_ni ix4974 (.Y (nx4973), .A0 (camera_module_cache_ram_216__1), .A1 (
             nx35180), .S0 (nx34522)) ;
    aoi22 ix29472 (.Y (nx29471), .A0 (camera_module_cache_ram_232__1), .A1 (
          nx36388), .B0 (camera_module_cache_ram_248__1), .B1 (nx36428)) ;
    dffr camera_module_cache_reg_ram_232__1 (.Q (camera_module_cache_ram_232__1)
         , .QB (\$dummy [1196]), .D (nx4963), .CLK (clk), .R (rst)) ;
    mux21_ni ix4964 (.Y (nx4963), .A0 (camera_module_cache_ram_232__1), .A1 (
             nx35180), .S0 (nx34518)) ;
    dffr camera_module_cache_reg_ram_248__1 (.Q (camera_module_cache_ram_248__1)
         , .QB (\$dummy [1197]), .D (nx4953), .CLK (clk), .R (rst)) ;
    mux21_ni ix4954 (.Y (nx4953), .A0 (camera_module_cache_ram_248__1), .A1 (
             nx35180), .S0 (nx34514)) ;
    oai21 ix29480 (.Y (nx29479), .A0 (nx7236), .A1 (nx7158), .B0 (nx36484)) ;
    nand04 ix7237 (.Y (nx7236), .A0 (nx29482), .A1 (nx29490), .A2 (nx29498), .A3 (
           nx29506)) ;
    aoi22 ix29483 (.Y (nx29482), .A0 (camera_module_cache_ram_9__1), .A1 (
          nx35830), .B0 (camera_module_cache_ram_25__1), .B1 (nx35870)) ;
    dffr camera_module_cache_reg_ram_9__1 (.Q (camera_module_cache_ram_9__1), .QB (
         \$dummy [1198]), .D (nx4943), .CLK (clk), .R (rst)) ;
    mux21_ni ix4944 (.Y (nx4943), .A0 (camera_module_cache_ram_9__1), .A1 (
             nx35180), .S0 (nx34504)) ;
    dffr camera_module_cache_reg_ram_25__1 (.Q (camera_module_cache_ram_25__1), 
         .QB (\$dummy [1199]), .D (nx4933), .CLK (clk), .R (rst)) ;
    mux21_ni ix4934 (.Y (nx4933), .A0 (camera_module_cache_ram_25__1), .A1 (
             nx35180), .S0 (nx34500)) ;
    aoi22 ix29491 (.Y (nx29490), .A0 (camera_module_cache_ram_41__1), .A1 (
          nx35910), .B0 (camera_module_cache_ram_57__1), .B1 (nx35950)) ;
    dffr camera_module_cache_reg_ram_41__1 (.Q (camera_module_cache_ram_41__1), 
         .QB (\$dummy [1200]), .D (nx4923), .CLK (clk), .R (rst)) ;
    mux21_ni ix4924 (.Y (nx4923), .A0 (camera_module_cache_ram_41__1), .A1 (
             nx35180), .S0 (nx34496)) ;
    dffr camera_module_cache_reg_ram_57__1 (.Q (camera_module_cache_ram_57__1), 
         .QB (\$dummy [1201]), .D (nx4913), .CLK (clk), .R (rst)) ;
    mux21_ni ix4914 (.Y (nx4913), .A0 (camera_module_cache_ram_57__1), .A1 (
             nx35182), .S0 (nx34492)) ;
    aoi22 ix29499 (.Y (nx29498), .A0 (camera_module_cache_ram_73__1), .A1 (
          nx35990), .B0 (camera_module_cache_ram_89__1), .B1 (nx36030)) ;
    dffr camera_module_cache_reg_ram_73__1 (.Q (camera_module_cache_ram_73__1), 
         .QB (\$dummy [1202]), .D (nx4903), .CLK (clk), .R (rst)) ;
    mux21_ni ix4904 (.Y (nx4903), .A0 (camera_module_cache_ram_73__1), .A1 (
             nx35182), .S0 (nx34488)) ;
    dffr camera_module_cache_reg_ram_89__1 (.Q (camera_module_cache_ram_89__1), 
         .QB (\$dummy [1203]), .D (nx4893), .CLK (clk), .R (rst)) ;
    mux21_ni ix4894 (.Y (nx4893), .A0 (camera_module_cache_ram_89__1), .A1 (
             nx35182), .S0 (nx34484)) ;
    aoi22 ix29507 (.Y (nx29506), .A0 (camera_module_cache_ram_121__1), .A1 (
          nx36070), .B0 (camera_module_cache_ram_105__1), .B1 (nx36110)) ;
    dffr camera_module_cache_reg_ram_121__1 (.Q (camera_module_cache_ram_121__1)
         , .QB (\$dummy [1204]), .D (nx4873), .CLK (clk), .R (rst)) ;
    mux21_ni ix4874 (.Y (nx4873), .A0 (camera_module_cache_ram_121__1), .A1 (
             nx35182), .S0 (nx34476)) ;
    dffr camera_module_cache_reg_ram_105__1 (.Q (camera_module_cache_ram_105__1)
         , .QB (\$dummy [1205]), .D (nx4883), .CLK (clk), .R (rst)) ;
    mux21_ni ix4884 (.Y (nx4883), .A0 (camera_module_cache_ram_105__1), .A1 (
             nx35182), .S0 (nx34480)) ;
    nand04 ix7159 (.Y (nx7158), .A0 (nx29515), .A1 (nx29523), .A2 (nx29531), .A3 (
           nx29539)) ;
    aoi22 ix29516 (.Y (nx29515), .A0 (camera_module_cache_ram_137__1), .A1 (
          nx36150), .B0 (camera_module_cache_ram_153__1), .B1 (nx36190)) ;
    dffr camera_module_cache_reg_ram_137__1 (.Q (camera_module_cache_ram_137__1)
         , .QB (\$dummy [1206]), .D (nx4863), .CLK (clk), .R (rst)) ;
    mux21_ni ix4864 (.Y (nx4863), .A0 (camera_module_cache_ram_137__1), .A1 (
             nx35182), .S0 (nx34472)) ;
    dffr camera_module_cache_reg_ram_153__1 (.Q (camera_module_cache_ram_153__1)
         , .QB (\$dummy [1207]), .D (nx4853), .CLK (clk), .R (rst)) ;
    mux21_ni ix4854 (.Y (nx4853), .A0 (camera_module_cache_ram_153__1), .A1 (
             nx35182), .S0 (nx34468)) ;
    aoi22 ix29524 (.Y (nx29523), .A0 (camera_module_cache_ram_185__1), .A1 (
          nx36230), .B0 (camera_module_cache_ram_169__1), .B1 (nx36270)) ;
    dffr camera_module_cache_reg_ram_185__1 (.Q (camera_module_cache_ram_185__1)
         , .QB (\$dummy [1208]), .D (nx4833), .CLK (clk), .R (rst)) ;
    mux21_ni ix4834 (.Y (nx4833), .A0 (camera_module_cache_ram_185__1), .A1 (
             nx35184), .S0 (nx34460)) ;
    dffr camera_module_cache_reg_ram_169__1 (.Q (camera_module_cache_ram_169__1)
         , .QB (\$dummy [1209]), .D (nx4843), .CLK (clk), .R (rst)) ;
    mux21_ni ix4844 (.Y (nx4843), .A0 (camera_module_cache_ram_169__1), .A1 (
             nx35184), .S0 (nx34464)) ;
    aoi22 ix29532 (.Y (nx29531), .A0 (camera_module_cache_ram_201__1), .A1 (
          nx36310), .B0 (camera_module_cache_ram_217__1), .B1 (nx36350)) ;
    dffr camera_module_cache_reg_ram_201__1 (.Q (camera_module_cache_ram_201__1)
         , .QB (\$dummy [1210]), .D (nx4823), .CLK (clk), .R (rst)) ;
    mux21_ni ix4824 (.Y (nx4823), .A0 (camera_module_cache_ram_201__1), .A1 (
             nx35184), .S0 (nx34456)) ;
    dffr camera_module_cache_reg_ram_217__1 (.Q (camera_module_cache_ram_217__1)
         , .QB (\$dummy [1211]), .D (nx4813), .CLK (clk), .R (rst)) ;
    mux21_ni ix4814 (.Y (nx4813), .A0 (camera_module_cache_ram_217__1), .A1 (
             nx35184), .S0 (nx34452)) ;
    aoi22 ix29540 (.Y (nx29539), .A0 (camera_module_cache_ram_233__1), .A1 (
          nx36390), .B0 (camera_module_cache_ram_249__1), .B1 (nx36430)) ;
    dffr camera_module_cache_reg_ram_233__1 (.Q (camera_module_cache_ram_233__1)
         , .QB (\$dummy [1212]), .D (nx4803), .CLK (clk), .R (rst)) ;
    mux21_ni ix4804 (.Y (nx4803), .A0 (camera_module_cache_ram_233__1), .A1 (
             nx35184), .S0 (nx34448)) ;
    dffr camera_module_cache_reg_ram_249__1 (.Q (camera_module_cache_ram_249__1)
         , .QB (\$dummy [1213]), .D (nx4793), .CLK (clk), .R (rst)) ;
    mux21_ni ix4794 (.Y (nx4793), .A0 (camera_module_cache_ram_249__1), .A1 (
             nx35184), .S0 (nx34444)) ;
    oai21 ix29548 (.Y (nx29547), .A0 (nx7072), .A1 (nx6994), .B0 (nx36488)) ;
    nand04 ix7073 (.Y (nx7072), .A0 (nx29550), .A1 (nx29558), .A2 (nx29566), .A3 (
           nx29574)) ;
    aoi22 ix29551 (.Y (nx29550), .A0 (camera_module_cache_ram_10__1), .A1 (
          nx35830), .B0 (camera_module_cache_ram_26__1), .B1 (nx35870)) ;
    dffr camera_module_cache_reg_ram_10__1 (.Q (camera_module_cache_ram_10__1), 
         .QB (\$dummy [1214]), .D (nx4783), .CLK (clk), .R (rst)) ;
    mux21_ni ix4784 (.Y (nx4783), .A0 (camera_module_cache_ram_10__1), .A1 (
             nx35184), .S0 (nx34434)) ;
    dffr camera_module_cache_reg_ram_26__1 (.Q (camera_module_cache_ram_26__1), 
         .QB (\$dummy [1215]), .D (nx4773), .CLK (clk), .R (rst)) ;
    mux21_ni ix4774 (.Y (nx4773), .A0 (camera_module_cache_ram_26__1), .A1 (
             nx35186), .S0 (nx34430)) ;
    aoi22 ix29559 (.Y (nx29558), .A0 (camera_module_cache_ram_42__1), .A1 (
          nx35910), .B0 (camera_module_cache_ram_58__1), .B1 (nx35950)) ;
    dffr camera_module_cache_reg_ram_42__1 (.Q (camera_module_cache_ram_42__1), 
         .QB (\$dummy [1216]), .D (nx4763), .CLK (clk), .R (rst)) ;
    mux21_ni ix4764 (.Y (nx4763), .A0 (camera_module_cache_ram_42__1), .A1 (
             nx35186), .S0 (nx34426)) ;
    dffr camera_module_cache_reg_ram_58__1 (.Q (camera_module_cache_ram_58__1), 
         .QB (\$dummy [1217]), .D (nx4753), .CLK (clk), .R (rst)) ;
    mux21_ni ix4754 (.Y (nx4753), .A0 (camera_module_cache_ram_58__1), .A1 (
             nx35186), .S0 (nx34422)) ;
    aoi22 ix29567 (.Y (nx29566), .A0 (camera_module_cache_ram_74__1), .A1 (
          nx35990), .B0 (camera_module_cache_ram_90__1), .B1 (nx36030)) ;
    dffr camera_module_cache_reg_ram_74__1 (.Q (camera_module_cache_ram_74__1), 
         .QB (\$dummy [1218]), .D (nx4743), .CLK (clk), .R (rst)) ;
    mux21_ni ix4744 (.Y (nx4743), .A0 (camera_module_cache_ram_74__1), .A1 (
             nx35186), .S0 (nx34418)) ;
    dffr camera_module_cache_reg_ram_90__1 (.Q (camera_module_cache_ram_90__1), 
         .QB (\$dummy [1219]), .D (nx4733), .CLK (clk), .R (rst)) ;
    mux21_ni ix4734 (.Y (nx4733), .A0 (camera_module_cache_ram_90__1), .A1 (
             nx35186), .S0 (nx34414)) ;
    aoi22 ix29575 (.Y (nx29574), .A0 (camera_module_cache_ram_122__1), .A1 (
          nx36070), .B0 (camera_module_cache_ram_106__1), .B1 (nx36110)) ;
    dffr camera_module_cache_reg_ram_122__1 (.Q (camera_module_cache_ram_122__1)
         , .QB (\$dummy [1220]), .D (nx4713), .CLK (clk), .R (rst)) ;
    mux21_ni ix4714 (.Y (nx4713), .A0 (camera_module_cache_ram_122__1), .A1 (
             nx35186), .S0 (nx34406)) ;
    dffr camera_module_cache_reg_ram_106__1 (.Q (camera_module_cache_ram_106__1)
         , .QB (\$dummy [1221]), .D (nx4723), .CLK (clk), .R (rst)) ;
    mux21_ni ix4724 (.Y (nx4723), .A0 (camera_module_cache_ram_106__1), .A1 (
             nx35186), .S0 (nx34410)) ;
    nand04 ix6995 (.Y (nx6994), .A0 (nx29583), .A1 (nx29591), .A2 (nx29599), .A3 (
           nx29607)) ;
    aoi22 ix29584 (.Y (nx29583), .A0 (camera_module_cache_ram_138__1), .A1 (
          nx36150), .B0 (camera_module_cache_ram_154__1), .B1 (nx36190)) ;
    dffr camera_module_cache_reg_ram_138__1 (.Q (camera_module_cache_ram_138__1)
         , .QB (\$dummy [1222]), .D (nx4703), .CLK (clk), .R (rst)) ;
    mux21_ni ix4704 (.Y (nx4703), .A0 (camera_module_cache_ram_138__1), .A1 (
             nx35188), .S0 (nx34402)) ;
    dffr camera_module_cache_reg_ram_154__1 (.Q (camera_module_cache_ram_154__1)
         , .QB (\$dummy [1223]), .D (nx4693), .CLK (clk), .R (rst)) ;
    mux21_ni ix4694 (.Y (nx4693), .A0 (camera_module_cache_ram_154__1), .A1 (
             nx35188), .S0 (nx34398)) ;
    aoi22 ix29592 (.Y (nx29591), .A0 (camera_module_cache_ram_186__1), .A1 (
          nx36230), .B0 (camera_module_cache_ram_170__1), .B1 (nx36270)) ;
    dffr camera_module_cache_reg_ram_186__1 (.Q (camera_module_cache_ram_186__1)
         , .QB (\$dummy [1224]), .D (nx4673), .CLK (clk), .R (rst)) ;
    mux21_ni ix4674 (.Y (nx4673), .A0 (camera_module_cache_ram_186__1), .A1 (
             nx35188), .S0 (nx34390)) ;
    dffr camera_module_cache_reg_ram_170__1 (.Q (camera_module_cache_ram_170__1)
         , .QB (\$dummy [1225]), .D (nx4683), .CLK (clk), .R (rst)) ;
    mux21_ni ix4684 (.Y (nx4683), .A0 (camera_module_cache_ram_170__1), .A1 (
             nx35188), .S0 (nx34394)) ;
    aoi22 ix29600 (.Y (nx29599), .A0 (camera_module_cache_ram_202__1), .A1 (
          nx36310), .B0 (camera_module_cache_ram_218__1), .B1 (nx36350)) ;
    dffr camera_module_cache_reg_ram_202__1 (.Q (camera_module_cache_ram_202__1)
         , .QB (\$dummy [1226]), .D (nx4663), .CLK (clk), .R (rst)) ;
    mux21_ni ix4664 (.Y (nx4663), .A0 (camera_module_cache_ram_202__1), .A1 (
             nx35188), .S0 (nx34386)) ;
    dffr camera_module_cache_reg_ram_218__1 (.Q (camera_module_cache_ram_218__1)
         , .QB (\$dummy [1227]), .D (nx4653), .CLK (clk), .R (rst)) ;
    mux21_ni ix4654 (.Y (nx4653), .A0 (camera_module_cache_ram_218__1), .A1 (
             nx35188), .S0 (nx34382)) ;
    aoi22 ix29608 (.Y (nx29607), .A0 (camera_module_cache_ram_234__1), .A1 (
          nx36390), .B0 (camera_module_cache_ram_250__1), .B1 (nx36430)) ;
    dffr camera_module_cache_reg_ram_234__1 (.Q (camera_module_cache_ram_234__1)
         , .QB (\$dummy [1228]), .D (nx4643), .CLK (clk), .R (rst)) ;
    mux21_ni ix4644 (.Y (nx4643), .A0 (camera_module_cache_ram_234__1), .A1 (
             nx35188), .S0 (nx34378)) ;
    dffr camera_module_cache_reg_ram_250__1 (.Q (camera_module_cache_ram_250__1)
         , .QB (\$dummy [1229]), .D (nx4633), .CLK (clk), .R (rst)) ;
    mux21_ni ix4634 (.Y (nx4633), .A0 (camera_module_cache_ram_250__1), .A1 (
             nx35190), .S0 (nx34374)) ;
    oai21 ix29616 (.Y (nx29615), .A0 (nx6910), .A1 (nx6832), .B0 (nx36492)) ;
    nand04 ix6911 (.Y (nx6910), .A0 (nx29618), .A1 (nx29626), .A2 (nx29634), .A3 (
           nx29642)) ;
    aoi22 ix29619 (.Y (nx29618), .A0 (camera_module_cache_ram_11__1), .A1 (
          nx35830), .B0 (camera_module_cache_ram_27__1), .B1 (nx35870)) ;
    dffr camera_module_cache_reg_ram_11__1 (.Q (camera_module_cache_ram_11__1), 
         .QB (\$dummy [1230]), .D (nx4623), .CLK (clk), .R (rst)) ;
    mux21_ni ix4624 (.Y (nx4623), .A0 (camera_module_cache_ram_11__1), .A1 (
             nx35190), .S0 (nx34364)) ;
    dffr camera_module_cache_reg_ram_27__1 (.Q (camera_module_cache_ram_27__1), 
         .QB (\$dummy [1231]), .D (nx4613), .CLK (clk), .R (rst)) ;
    mux21_ni ix4614 (.Y (nx4613), .A0 (camera_module_cache_ram_27__1), .A1 (
             nx35190), .S0 (nx34360)) ;
    aoi22 ix29627 (.Y (nx29626), .A0 (camera_module_cache_ram_43__1), .A1 (
          nx35910), .B0 (camera_module_cache_ram_59__1), .B1 (nx35950)) ;
    dffr camera_module_cache_reg_ram_43__1 (.Q (camera_module_cache_ram_43__1), 
         .QB (\$dummy [1232]), .D (nx4603), .CLK (clk), .R (rst)) ;
    mux21_ni ix4604 (.Y (nx4603), .A0 (camera_module_cache_ram_43__1), .A1 (
             nx35190), .S0 (nx34356)) ;
    dffr camera_module_cache_reg_ram_59__1 (.Q (camera_module_cache_ram_59__1), 
         .QB (\$dummy [1233]), .D (nx4593), .CLK (clk), .R (rst)) ;
    mux21_ni ix4594 (.Y (nx4593), .A0 (camera_module_cache_ram_59__1), .A1 (
             nx35190), .S0 (nx34352)) ;
    aoi22 ix29635 (.Y (nx29634), .A0 (camera_module_cache_ram_75__1), .A1 (
          nx35990), .B0 (camera_module_cache_ram_91__1), .B1 (nx36030)) ;
    dffr camera_module_cache_reg_ram_75__1 (.Q (camera_module_cache_ram_75__1), 
         .QB (\$dummy [1234]), .D (nx4583), .CLK (clk), .R (rst)) ;
    mux21_ni ix4584 (.Y (nx4583), .A0 (camera_module_cache_ram_75__1), .A1 (
             nx35190), .S0 (nx34348)) ;
    dffr camera_module_cache_reg_ram_91__1 (.Q (camera_module_cache_ram_91__1), 
         .QB (\$dummy [1235]), .D (nx4573), .CLK (clk), .R (rst)) ;
    mux21_ni ix4574 (.Y (nx4573), .A0 (camera_module_cache_ram_91__1), .A1 (
             nx35190), .S0 (nx34344)) ;
    aoi22 ix29643 (.Y (nx29642), .A0 (camera_module_cache_ram_123__1), .A1 (
          nx36070), .B0 (camera_module_cache_ram_107__1), .B1 (nx36110)) ;
    dffr camera_module_cache_reg_ram_123__1 (.Q (camera_module_cache_ram_123__1)
         , .QB (\$dummy [1236]), .D (nx4553), .CLK (clk), .R (rst)) ;
    mux21_ni ix4554 (.Y (nx4553), .A0 (camera_module_cache_ram_123__1), .A1 (
             nx35192), .S0 (nx34336)) ;
    dffr camera_module_cache_reg_ram_107__1 (.Q (camera_module_cache_ram_107__1)
         , .QB (\$dummy [1237]), .D (nx4563), .CLK (clk), .R (rst)) ;
    mux21_ni ix4564 (.Y (nx4563), .A0 (camera_module_cache_ram_107__1), .A1 (
             nx35192), .S0 (nx34340)) ;
    nand04 ix6833 (.Y (nx6832), .A0 (nx29651), .A1 (nx29659), .A2 (nx29667), .A3 (
           nx29675)) ;
    aoi22 ix29652 (.Y (nx29651), .A0 (camera_module_cache_ram_139__1), .A1 (
          nx36150), .B0 (camera_module_cache_ram_155__1), .B1 (nx36190)) ;
    dffr camera_module_cache_reg_ram_139__1 (.Q (camera_module_cache_ram_139__1)
         , .QB (\$dummy [1238]), .D (nx4543), .CLK (clk), .R (rst)) ;
    mux21_ni ix4544 (.Y (nx4543), .A0 (camera_module_cache_ram_139__1), .A1 (
             nx35192), .S0 (nx34332)) ;
    dffr camera_module_cache_reg_ram_155__1 (.Q (camera_module_cache_ram_155__1)
         , .QB (\$dummy [1239]), .D (nx4533), .CLK (clk), .R (rst)) ;
    mux21_ni ix4534 (.Y (nx4533), .A0 (camera_module_cache_ram_155__1), .A1 (
             nx35192), .S0 (nx34328)) ;
    aoi22 ix29660 (.Y (nx29659), .A0 (camera_module_cache_ram_187__1), .A1 (
          nx36230), .B0 (camera_module_cache_ram_171__1), .B1 (nx36270)) ;
    dffr camera_module_cache_reg_ram_187__1 (.Q (camera_module_cache_ram_187__1)
         , .QB (\$dummy [1240]), .D (nx4513), .CLK (clk), .R (rst)) ;
    mux21_ni ix4514 (.Y (nx4513), .A0 (camera_module_cache_ram_187__1), .A1 (
             nx35192), .S0 (nx34320)) ;
    dffr camera_module_cache_reg_ram_171__1 (.Q (camera_module_cache_ram_171__1)
         , .QB (\$dummy [1241]), .D (nx4523), .CLK (clk), .R (rst)) ;
    mux21_ni ix4524 (.Y (nx4523), .A0 (camera_module_cache_ram_171__1), .A1 (
             nx35192), .S0 (nx34324)) ;
    aoi22 ix29668 (.Y (nx29667), .A0 (camera_module_cache_ram_203__1), .A1 (
          nx36310), .B0 (camera_module_cache_ram_219__1), .B1 (nx36350)) ;
    dffr camera_module_cache_reg_ram_203__1 (.Q (camera_module_cache_ram_203__1)
         , .QB (\$dummy [1242]), .D (nx4503), .CLK (clk), .R (rst)) ;
    mux21_ni ix4504 (.Y (nx4503), .A0 (camera_module_cache_ram_203__1), .A1 (
             nx35192), .S0 (nx34316)) ;
    dffr camera_module_cache_reg_ram_219__1 (.Q (camera_module_cache_ram_219__1)
         , .QB (\$dummy [1243]), .D (nx4493), .CLK (clk), .R (rst)) ;
    mux21_ni ix4494 (.Y (nx4493), .A0 (camera_module_cache_ram_219__1), .A1 (
             nx35194), .S0 (nx34312)) ;
    aoi22 ix29676 (.Y (nx29675), .A0 (camera_module_cache_ram_235__1), .A1 (
          nx36390), .B0 (camera_module_cache_ram_251__1), .B1 (nx36430)) ;
    dffr camera_module_cache_reg_ram_235__1 (.Q (camera_module_cache_ram_235__1)
         , .QB (\$dummy [1244]), .D (nx4483), .CLK (clk), .R (rst)) ;
    mux21_ni ix4484 (.Y (nx4483), .A0 (camera_module_cache_ram_235__1), .A1 (
             nx35194), .S0 (nx34308)) ;
    dffr camera_module_cache_reg_ram_251__1 (.Q (camera_module_cache_ram_251__1)
         , .QB (\$dummy [1245]), .D (nx4473), .CLK (clk), .R (rst)) ;
    mux21_ni ix4474 (.Y (nx4473), .A0 (camera_module_cache_ram_251__1), .A1 (
             nx35194), .S0 (nx34304)) ;
    nand04 ix6755 (.Y (nx6754), .A0 (nx29684), .A1 (nx29752), .A2 (nx29820), .A3 (
           nx29888)) ;
    oai21 ix29685 (.Y (nx29684), .A0 (nx6744), .A1 (nx6666), .B0 (nx36506)) ;
    nand04 ix6745 (.Y (nx6744), .A0 (nx29687), .A1 (nx29695), .A2 (nx29703), .A3 (
           nx29711)) ;
    aoi22 ix29688 (.Y (nx29687), .A0 (camera_module_cache_ram_12__1), .A1 (
          nx35830), .B0 (camera_module_cache_ram_28__1), .B1 (nx35870)) ;
    dffr camera_module_cache_reg_ram_12__1 (.Q (camera_module_cache_ram_12__1), 
         .QB (\$dummy [1246]), .D (nx4463), .CLK (clk), .R (rst)) ;
    mux21_ni ix4464 (.Y (nx4463), .A0 (nx35194), .A1 (
             camera_module_cache_ram_12__1), .S0 (nx36496)) ;
    dffr camera_module_cache_reg_ram_28__1 (.Q (camera_module_cache_ram_28__1), 
         .QB (\$dummy [1247]), .D (nx4453), .CLK (clk), .R (rst)) ;
    mux21_ni ix4454 (.Y (nx4453), .A0 (nx35194), .A1 (
             camera_module_cache_ram_28__1), .S0 (nx36510)) ;
    aoi22 ix29696 (.Y (nx29695), .A0 (camera_module_cache_ram_44__1), .A1 (
          nx35910), .B0 (camera_module_cache_ram_60__1), .B1 (nx35950)) ;
    dffr camera_module_cache_reg_ram_44__1 (.Q (camera_module_cache_ram_44__1), 
         .QB (\$dummy [1248]), .D (nx4443), .CLK (clk), .R (rst)) ;
    mux21_ni ix4444 (.Y (nx4443), .A0 (nx35194), .A1 (
             camera_module_cache_ram_44__1), .S0 (nx36514)) ;
    dffr camera_module_cache_reg_ram_60__1 (.Q (camera_module_cache_ram_60__1), 
         .QB (\$dummy [1249]), .D (nx4433), .CLK (clk), .R (rst)) ;
    mux21_ni ix4434 (.Y (nx4433), .A0 (nx35194), .A1 (
             camera_module_cache_ram_60__1), .S0 (nx36518)) ;
    aoi22 ix29704 (.Y (nx29703), .A0 (camera_module_cache_ram_76__1), .A1 (
          nx35990), .B0 (camera_module_cache_ram_92__1), .B1 (nx36030)) ;
    dffr camera_module_cache_reg_ram_76__1 (.Q (camera_module_cache_ram_76__1), 
         .QB (\$dummy [1250]), .D (nx4423), .CLK (clk), .R (rst)) ;
    mux21_ni ix4424 (.Y (nx4423), .A0 (nx35196), .A1 (
             camera_module_cache_ram_76__1), .S0 (nx36522)) ;
    dffr camera_module_cache_reg_ram_92__1 (.Q (camera_module_cache_ram_92__1), 
         .QB (\$dummy [1251]), .D (nx4413), .CLK (clk), .R (rst)) ;
    mux21_ni ix4414 (.Y (nx4413), .A0 (nx35196), .A1 (
             camera_module_cache_ram_92__1), .S0 (nx36526)) ;
    aoi22 ix29712 (.Y (nx29711), .A0 (camera_module_cache_ram_124__1), .A1 (
          nx36070), .B0 (camera_module_cache_ram_108__1), .B1 (nx36110)) ;
    dffr camera_module_cache_reg_ram_124__1 (.Q (camera_module_cache_ram_124__1)
         , .QB (\$dummy [1252]), .D (nx4393), .CLK (clk), .R (rst)) ;
    mux21_ni ix4394 (.Y (nx4393), .A0 (nx35196), .A1 (
             camera_module_cache_ram_124__1), .S0 (nx36530)) ;
    dffr camera_module_cache_reg_ram_108__1 (.Q (camera_module_cache_ram_108__1)
         , .QB (\$dummy [1253]), .D (nx4403), .CLK (clk), .R (rst)) ;
    mux21_ni ix4404 (.Y (nx4403), .A0 (nx35196), .A1 (
             camera_module_cache_ram_108__1), .S0 (nx36534)) ;
    nand04 ix6667 (.Y (nx6666), .A0 (nx29720), .A1 (nx29728), .A2 (nx29736), .A3 (
           nx29744)) ;
    aoi22 ix29721 (.Y (nx29720), .A0 (camera_module_cache_ram_140__1), .A1 (
          nx36150), .B0 (camera_module_cache_ram_156__1), .B1 (nx36190)) ;
    dffr camera_module_cache_reg_ram_140__1 (.Q (camera_module_cache_ram_140__1)
         , .QB (\$dummy [1254]), .D (nx4383), .CLK (clk), .R (rst)) ;
    mux21_ni ix4384 (.Y (nx4383), .A0 (nx35196), .A1 (
             camera_module_cache_ram_140__1), .S0 (nx36538)) ;
    dffr camera_module_cache_reg_ram_156__1 (.Q (camera_module_cache_ram_156__1)
         , .QB (\$dummy [1255]), .D (nx4373), .CLK (clk), .R (rst)) ;
    mux21_ni ix4374 (.Y (nx4373), .A0 (nx35196), .A1 (
             camera_module_cache_ram_156__1), .S0 (nx36542)) ;
    aoi22 ix29729 (.Y (nx29728), .A0 (camera_module_cache_ram_188__1), .A1 (
          nx36230), .B0 (camera_module_cache_ram_172__1), .B1 (nx36270)) ;
    dffr camera_module_cache_reg_ram_188__1 (.Q (camera_module_cache_ram_188__1)
         , .QB (\$dummy [1256]), .D (nx4353), .CLK (clk), .R (rst)) ;
    mux21_ni ix4354 (.Y (nx4353), .A0 (nx35196), .A1 (
             camera_module_cache_ram_188__1), .S0 (nx36546)) ;
    dffr camera_module_cache_reg_ram_172__1 (.Q (camera_module_cache_ram_172__1)
         , .QB (\$dummy [1257]), .D (nx4363), .CLK (clk), .R (rst)) ;
    mux21_ni ix4364 (.Y (nx4363), .A0 (nx35198), .A1 (
             camera_module_cache_ram_172__1), .S0 (nx36550)) ;
    aoi22 ix29737 (.Y (nx29736), .A0 (camera_module_cache_ram_204__1), .A1 (
          nx36310), .B0 (camera_module_cache_ram_220__1), .B1 (nx36350)) ;
    dffr camera_module_cache_reg_ram_204__1 (.Q (camera_module_cache_ram_204__1)
         , .QB (\$dummy [1258]), .D (nx4343), .CLK (clk), .R (rst)) ;
    mux21_ni ix4344 (.Y (nx4343), .A0 (nx35198), .A1 (
             camera_module_cache_ram_204__1), .S0 (nx36554)) ;
    dffr camera_module_cache_reg_ram_220__1 (.Q (camera_module_cache_ram_220__1)
         , .QB (\$dummy [1259]), .D (nx4333), .CLK (clk), .R (rst)) ;
    mux21_ni ix4334 (.Y (nx4333), .A0 (nx35198), .A1 (
             camera_module_cache_ram_220__1), .S0 (nx36558)) ;
    aoi22 ix29745 (.Y (nx29744), .A0 (camera_module_cache_ram_236__1), .A1 (
          nx36390), .B0 (camera_module_cache_ram_252__1), .B1 (nx36430)) ;
    dffr camera_module_cache_reg_ram_236__1 (.Q (camera_module_cache_ram_236__1)
         , .QB (\$dummy [1260]), .D (nx4323), .CLK (clk), .R (rst)) ;
    mux21_ni ix4324 (.Y (nx4323), .A0 (nx35198), .A1 (
             camera_module_cache_ram_236__1), .S0 (nx36562)) ;
    dffr camera_module_cache_reg_ram_252__1 (.Q (camera_module_cache_ram_252__1)
         , .QB (\$dummy [1261]), .D (nx4313), .CLK (clk), .R (rst)) ;
    mux21_ni ix4314 (.Y (nx4313), .A0 (nx35198), .A1 (
             camera_module_cache_ram_252__1), .S0 (nx36566)) ;
    oai21 ix29753 (.Y (nx29752), .A0 (nx6582), .A1 (nx6504), .B0 (nx36580)) ;
    nand04 ix6583 (.Y (nx6582), .A0 (nx29755), .A1 (nx29763), .A2 (nx29771), .A3 (
           nx29779)) ;
    aoi22 ix29756 (.Y (nx29755), .A0 (camera_module_cache_ram_13__1), .A1 (
          nx35830), .B0 (camera_module_cache_ram_29__1), .B1 (nx35870)) ;
    dffr camera_module_cache_reg_ram_13__1 (.Q (camera_module_cache_ram_13__1), 
         .QB (\$dummy [1262]), .D (nx4303), .CLK (clk), .R (rst)) ;
    mux21_ni ix4304 (.Y (nx4303), .A0 (nx35198), .A1 (
             camera_module_cache_ram_13__1), .S0 (nx36570)) ;
    dffr camera_module_cache_reg_ram_29__1 (.Q (camera_module_cache_ram_29__1), 
         .QB (\$dummy [1263]), .D (nx4293), .CLK (clk), .R (rst)) ;
    mux21_ni ix4294 (.Y (nx4293), .A0 (nx35198), .A1 (
             camera_module_cache_ram_29__1), .S0 (nx36584)) ;
    aoi22 ix29764 (.Y (nx29763), .A0 (camera_module_cache_ram_45__1), .A1 (
          nx35910), .B0 (camera_module_cache_ram_61__1), .B1 (nx35950)) ;
    dffr camera_module_cache_reg_ram_45__1 (.Q (camera_module_cache_ram_45__1), 
         .QB (\$dummy [1264]), .D (nx4283), .CLK (clk), .R (rst)) ;
    mux21_ni ix4284 (.Y (nx4283), .A0 (nx35200), .A1 (
             camera_module_cache_ram_45__1), .S0 (nx36588)) ;
    dffr camera_module_cache_reg_ram_61__1 (.Q (camera_module_cache_ram_61__1), 
         .QB (\$dummy [1265]), .D (nx4273), .CLK (clk), .R (rst)) ;
    mux21_ni ix4274 (.Y (nx4273), .A0 (nx35200), .A1 (
             camera_module_cache_ram_61__1), .S0 (nx36592)) ;
    aoi22 ix29772 (.Y (nx29771), .A0 (camera_module_cache_ram_77__1), .A1 (
          nx35990), .B0 (camera_module_cache_ram_93__1), .B1 (nx36030)) ;
    dffr camera_module_cache_reg_ram_77__1 (.Q (camera_module_cache_ram_77__1), 
         .QB (\$dummy [1266]), .D (nx4263), .CLK (clk), .R (rst)) ;
    mux21_ni ix4264 (.Y (nx4263), .A0 (nx35200), .A1 (
             camera_module_cache_ram_77__1), .S0 (nx36596)) ;
    dffr camera_module_cache_reg_ram_93__1 (.Q (camera_module_cache_ram_93__1), 
         .QB (\$dummy [1267]), .D (nx4253), .CLK (clk), .R (rst)) ;
    mux21_ni ix4254 (.Y (nx4253), .A0 (nx35200), .A1 (
             camera_module_cache_ram_93__1), .S0 (nx36600)) ;
    aoi22 ix29780 (.Y (nx29779), .A0 (camera_module_cache_ram_125__1), .A1 (
          nx36070), .B0 (camera_module_cache_ram_109__1), .B1 (nx36110)) ;
    dffr camera_module_cache_reg_ram_125__1 (.Q (camera_module_cache_ram_125__1)
         , .QB (\$dummy [1268]), .D (nx4233), .CLK (clk), .R (rst)) ;
    mux21_ni ix4234 (.Y (nx4233), .A0 (nx35200), .A1 (
             camera_module_cache_ram_125__1), .S0 (nx36604)) ;
    dffr camera_module_cache_reg_ram_109__1 (.Q (camera_module_cache_ram_109__1)
         , .QB (\$dummy [1269]), .D (nx4243), .CLK (clk), .R (rst)) ;
    mux21_ni ix4244 (.Y (nx4243), .A0 (nx35200), .A1 (
             camera_module_cache_ram_109__1), .S0 (nx36608)) ;
    nand04 ix6505 (.Y (nx6504), .A0 (nx29788), .A1 (nx29796), .A2 (nx29804), .A3 (
           nx29812)) ;
    aoi22 ix29789 (.Y (nx29788), .A0 (camera_module_cache_ram_141__1), .A1 (
          nx36150), .B0 (camera_module_cache_ram_157__1), .B1 (nx36190)) ;
    dffr camera_module_cache_reg_ram_141__1 (.Q (camera_module_cache_ram_141__1)
         , .QB (\$dummy [1270]), .D (nx4223), .CLK (clk), .R (rst)) ;
    mux21_ni ix4224 (.Y (nx4223), .A0 (nx35200), .A1 (
             camera_module_cache_ram_141__1), .S0 (nx36612)) ;
    dffr camera_module_cache_reg_ram_157__1 (.Q (camera_module_cache_ram_157__1)
         , .QB (\$dummy [1271]), .D (nx4213), .CLK (clk), .R (rst)) ;
    mux21_ni ix4214 (.Y (nx4213), .A0 (nx35202), .A1 (
             camera_module_cache_ram_157__1), .S0 (nx36616)) ;
    aoi22 ix29797 (.Y (nx29796), .A0 (camera_module_cache_ram_189__1), .A1 (
          nx36230), .B0 (camera_module_cache_ram_173__1), .B1 (nx36270)) ;
    dffr camera_module_cache_reg_ram_189__1 (.Q (camera_module_cache_ram_189__1)
         , .QB (\$dummy [1272]), .D (nx4193), .CLK (clk), .R (rst)) ;
    mux21_ni ix4194 (.Y (nx4193), .A0 (nx35202), .A1 (
             camera_module_cache_ram_189__1), .S0 (nx36620)) ;
    dffr camera_module_cache_reg_ram_173__1 (.Q (camera_module_cache_ram_173__1)
         , .QB (\$dummy [1273]), .D (nx4203), .CLK (clk), .R (rst)) ;
    mux21_ni ix4204 (.Y (nx4203), .A0 (nx35202), .A1 (
             camera_module_cache_ram_173__1), .S0 (nx36624)) ;
    aoi22 ix29805 (.Y (nx29804), .A0 (camera_module_cache_ram_205__1), .A1 (
          nx36310), .B0 (camera_module_cache_ram_221__1), .B1 (nx36350)) ;
    dffr camera_module_cache_reg_ram_205__1 (.Q (camera_module_cache_ram_205__1)
         , .QB (\$dummy [1274]), .D (nx4183), .CLK (clk), .R (rst)) ;
    mux21_ni ix4184 (.Y (nx4183), .A0 (nx35202), .A1 (
             camera_module_cache_ram_205__1), .S0 (nx36628)) ;
    dffr camera_module_cache_reg_ram_221__1 (.Q (camera_module_cache_ram_221__1)
         , .QB (\$dummy [1275]), .D (nx4173), .CLK (clk), .R (rst)) ;
    mux21_ni ix4174 (.Y (nx4173), .A0 (nx35202), .A1 (
             camera_module_cache_ram_221__1), .S0 (nx36632)) ;
    aoi22 ix29813 (.Y (nx29812), .A0 (camera_module_cache_ram_237__1), .A1 (
          nx36390), .B0 (camera_module_cache_ram_253__1), .B1 (nx36430)) ;
    dffr camera_module_cache_reg_ram_237__1 (.Q (camera_module_cache_ram_237__1)
         , .QB (\$dummy [1276]), .D (nx4163), .CLK (clk), .R (rst)) ;
    mux21_ni ix4164 (.Y (nx4163), .A0 (nx35202), .A1 (
             camera_module_cache_ram_237__1), .S0 (nx36636)) ;
    dffr camera_module_cache_reg_ram_253__1 (.Q (camera_module_cache_ram_253__1)
         , .QB (\$dummy [1277]), .D (nx4153), .CLK (clk), .R (rst)) ;
    mux21_ni ix4154 (.Y (nx4153), .A0 (nx35202), .A1 (
             camera_module_cache_ram_253__1), .S0 (nx36640)) ;
    oai21 ix29821 (.Y (nx29820), .A0 (nx6418), .A1 (nx6340), .B0 (nx36654)) ;
    nand04 ix6419 (.Y (nx6418), .A0 (nx29823), .A1 (nx29831), .A2 (nx29839), .A3 (
           nx29847)) ;
    aoi22 ix29824 (.Y (nx29823), .A0 (camera_module_cache_ram_14__1), .A1 (
          nx35830), .B0 (camera_module_cache_ram_30__1), .B1 (nx35870)) ;
    dffr camera_module_cache_reg_ram_14__1 (.Q (camera_module_cache_ram_14__1), 
         .QB (\$dummy [1278]), .D (nx4143), .CLK (clk), .R (rst)) ;
    mux21_ni ix4144 (.Y (nx4143), .A0 (nx35204), .A1 (
             camera_module_cache_ram_14__1), .S0 (nx36644)) ;
    dffr camera_module_cache_reg_ram_30__1 (.Q (camera_module_cache_ram_30__1), 
         .QB (\$dummy [1279]), .D (nx4133), .CLK (clk), .R (rst)) ;
    mux21_ni ix4134 (.Y (nx4133), .A0 (nx35204), .A1 (
             camera_module_cache_ram_30__1), .S0 (nx36658)) ;
    aoi22 ix29832 (.Y (nx29831), .A0 (camera_module_cache_ram_46__1), .A1 (
          nx35910), .B0 (camera_module_cache_ram_62__1), .B1 (nx35950)) ;
    dffr camera_module_cache_reg_ram_46__1 (.Q (camera_module_cache_ram_46__1), 
         .QB (\$dummy [1280]), .D (nx4123), .CLK (clk), .R (rst)) ;
    mux21_ni ix4124 (.Y (nx4123), .A0 (nx35204), .A1 (
             camera_module_cache_ram_46__1), .S0 (nx36662)) ;
    dffr camera_module_cache_reg_ram_62__1 (.Q (camera_module_cache_ram_62__1), 
         .QB (\$dummy [1281]), .D (nx4113), .CLK (clk), .R (rst)) ;
    mux21_ni ix4114 (.Y (nx4113), .A0 (nx35204), .A1 (
             camera_module_cache_ram_62__1), .S0 (nx36666)) ;
    aoi22 ix29840 (.Y (nx29839), .A0 (camera_module_cache_ram_78__1), .A1 (
          nx35990), .B0 (camera_module_cache_ram_94__1), .B1 (nx36030)) ;
    dffr camera_module_cache_reg_ram_78__1 (.Q (camera_module_cache_ram_78__1), 
         .QB (\$dummy [1282]), .D (nx4103), .CLK (clk), .R (rst)) ;
    mux21_ni ix4104 (.Y (nx4103), .A0 (nx35204), .A1 (
             camera_module_cache_ram_78__1), .S0 (nx36670)) ;
    dffr camera_module_cache_reg_ram_94__1 (.Q (camera_module_cache_ram_94__1), 
         .QB (\$dummy [1283]), .D (nx4093), .CLK (clk), .R (rst)) ;
    mux21_ni ix4094 (.Y (nx4093), .A0 (nx35204), .A1 (
             camera_module_cache_ram_94__1), .S0 (nx36674)) ;
    aoi22 ix29848 (.Y (nx29847), .A0 (camera_module_cache_ram_126__1), .A1 (
          nx36070), .B0 (camera_module_cache_ram_110__1), .B1 (nx36110)) ;
    dffr camera_module_cache_reg_ram_126__1 (.Q (camera_module_cache_ram_126__1)
         , .QB (\$dummy [1284]), .D (nx4073), .CLK (clk), .R (rst)) ;
    mux21_ni ix4074 (.Y (nx4073), .A0 (nx35204), .A1 (
             camera_module_cache_ram_126__1), .S0 (nx36678)) ;
    dffr camera_module_cache_reg_ram_110__1 (.Q (camera_module_cache_ram_110__1)
         , .QB (\$dummy [1285]), .D (nx4083), .CLK (clk), .R (rst)) ;
    mux21_ni ix4084 (.Y (nx4083), .A0 (nx35206), .A1 (
             camera_module_cache_ram_110__1), .S0 (nx36682)) ;
    nand04 ix6341 (.Y (nx6340), .A0 (nx29856), .A1 (nx29864), .A2 (nx29872), .A3 (
           nx29880)) ;
    aoi22 ix29857 (.Y (nx29856), .A0 (camera_module_cache_ram_142__1), .A1 (
          nx36150), .B0 (camera_module_cache_ram_158__1), .B1 (nx36190)) ;
    dffr camera_module_cache_reg_ram_142__1 (.Q (camera_module_cache_ram_142__1)
         , .QB (\$dummy [1286]), .D (nx4063), .CLK (clk), .R (rst)) ;
    mux21_ni ix4064 (.Y (nx4063), .A0 (nx35206), .A1 (
             camera_module_cache_ram_142__1), .S0 (nx36686)) ;
    dffr camera_module_cache_reg_ram_158__1 (.Q (camera_module_cache_ram_158__1)
         , .QB (\$dummy [1287]), .D (nx4053), .CLK (clk), .R (rst)) ;
    mux21_ni ix4054 (.Y (nx4053), .A0 (nx35206), .A1 (
             camera_module_cache_ram_158__1), .S0 (nx36690)) ;
    aoi22 ix29865 (.Y (nx29864), .A0 (camera_module_cache_ram_190__1), .A1 (
          nx36230), .B0 (camera_module_cache_ram_174__1), .B1 (nx36270)) ;
    dffr camera_module_cache_reg_ram_190__1 (.Q (camera_module_cache_ram_190__1)
         , .QB (\$dummy [1288]), .D (nx4033), .CLK (clk), .R (rst)) ;
    mux21_ni ix4034 (.Y (nx4033), .A0 (nx35206), .A1 (
             camera_module_cache_ram_190__1), .S0 (nx36694)) ;
    dffr camera_module_cache_reg_ram_174__1 (.Q (camera_module_cache_ram_174__1)
         , .QB (\$dummy [1289]), .D (nx4043), .CLK (clk), .R (rst)) ;
    mux21_ni ix4044 (.Y (nx4043), .A0 (nx35206), .A1 (
             camera_module_cache_ram_174__1), .S0 (nx36698)) ;
    aoi22 ix29873 (.Y (nx29872), .A0 (camera_module_cache_ram_206__1), .A1 (
          nx36310), .B0 (camera_module_cache_ram_222__1), .B1 (nx36350)) ;
    dffr camera_module_cache_reg_ram_206__1 (.Q (camera_module_cache_ram_206__1)
         , .QB (\$dummy [1290]), .D (nx4023), .CLK (clk), .R (rst)) ;
    mux21_ni ix4024 (.Y (nx4023), .A0 (nx35206), .A1 (
             camera_module_cache_ram_206__1), .S0 (nx36702)) ;
    dffr camera_module_cache_reg_ram_222__1 (.Q (camera_module_cache_ram_222__1)
         , .QB (\$dummy [1291]), .D (nx4013), .CLK (clk), .R (rst)) ;
    mux21_ni ix4014 (.Y (nx4013), .A0 (nx35206), .A1 (
             camera_module_cache_ram_222__1), .S0 (nx36706)) ;
    aoi22 ix29881 (.Y (nx29880), .A0 (camera_module_cache_ram_238__1), .A1 (
          nx36390), .B0 (camera_module_cache_ram_254__1), .B1 (nx36430)) ;
    dffr camera_module_cache_reg_ram_238__1 (.Q (camera_module_cache_ram_238__1)
         , .QB (\$dummy [1292]), .D (nx4003), .CLK (clk), .R (rst)) ;
    mux21_ni ix4004 (.Y (nx4003), .A0 (nx35208), .A1 (
             camera_module_cache_ram_238__1), .S0 (nx36710)) ;
    dffr camera_module_cache_reg_ram_254__1 (.Q (camera_module_cache_ram_254__1)
         , .QB (\$dummy [1293]), .D (nx3993), .CLK (clk), .R (rst)) ;
    mux21_ni ix3994 (.Y (nx3993), .A0 (nx35208), .A1 (
             camera_module_cache_ram_254__1), .S0 (nx36714)) ;
    oai21 ix29889 (.Y (nx29888), .A0 (nx6256), .A1 (nx6178), .B0 (nx36728)) ;
    nand04 ix6257 (.Y (nx6256), .A0 (nx29891), .A1 (nx29899), .A2 (nx29907), .A3 (
           nx29915)) ;
    aoi22 ix29892 (.Y (nx29891), .A0 (camera_module_cache_ram_15__1), .A1 (
          nx35830), .B0 (camera_module_cache_ram_31__1), .B1 (nx35870)) ;
    dffr camera_module_cache_reg_ram_15__1 (.Q (camera_module_cache_ram_15__1), 
         .QB (\$dummy [1294]), .D (nx3983), .CLK (clk), .R (rst)) ;
    mux21_ni ix3984 (.Y (nx3983), .A0 (nx35208), .A1 (
             camera_module_cache_ram_15__1), .S0 (nx36718)) ;
    dffr camera_module_cache_reg_ram_31__1 (.Q (camera_module_cache_ram_31__1), 
         .QB (\$dummy [1295]), .D (nx3973), .CLK (clk), .R (rst)) ;
    mux21_ni ix3974 (.Y (nx3973), .A0 (nx35208), .A1 (
             camera_module_cache_ram_31__1), .S0 (nx36732)) ;
    aoi22 ix29900 (.Y (nx29899), .A0 (camera_module_cache_ram_47__1), .A1 (
          nx35910), .B0 (camera_module_cache_ram_63__1), .B1 (nx35950)) ;
    dffr camera_module_cache_reg_ram_47__1 (.Q (camera_module_cache_ram_47__1), 
         .QB (\$dummy [1296]), .D (nx3963), .CLK (clk), .R (rst)) ;
    mux21_ni ix3964 (.Y (nx3963), .A0 (nx35208), .A1 (
             camera_module_cache_ram_47__1), .S0 (nx36736)) ;
    dffr camera_module_cache_reg_ram_63__1 (.Q (camera_module_cache_ram_63__1), 
         .QB (\$dummy [1297]), .D (nx3953), .CLK (clk), .R (rst)) ;
    mux21_ni ix3954 (.Y (nx3953), .A0 (nx35208), .A1 (
             camera_module_cache_ram_63__1), .S0 (nx36740)) ;
    aoi22 ix29908 (.Y (nx29907), .A0 (camera_module_cache_ram_79__1), .A1 (
          nx35990), .B0 (camera_module_cache_ram_95__1), .B1 (nx36030)) ;
    dffr camera_module_cache_reg_ram_79__1 (.Q (camera_module_cache_ram_79__1), 
         .QB (\$dummy [1298]), .D (nx3943), .CLK (clk), .R (rst)) ;
    mux21_ni ix3944 (.Y (nx3943), .A0 (nx35208), .A1 (
             camera_module_cache_ram_79__1), .S0 (nx36744)) ;
    dffr camera_module_cache_reg_ram_95__1 (.Q (camera_module_cache_ram_95__1), 
         .QB (\$dummy [1299]), .D (nx3933), .CLK (clk), .R (rst)) ;
    mux21_ni ix3934 (.Y (nx3933), .A0 (nx35210), .A1 (
             camera_module_cache_ram_95__1), .S0 (nx36748)) ;
    aoi22 ix29916 (.Y (nx29915), .A0 (camera_module_cache_ram_127__1), .A1 (
          nx36070), .B0 (camera_module_cache_ram_111__1), .B1 (nx36110)) ;
    dffr camera_module_cache_reg_ram_127__1 (.Q (camera_module_cache_ram_127__1)
         , .QB (\$dummy [1300]), .D (nx3913), .CLK (clk), .R (rst)) ;
    mux21_ni ix3914 (.Y (nx3913), .A0 (nx35210), .A1 (
             camera_module_cache_ram_127__1), .S0 (nx36752)) ;
    dffr camera_module_cache_reg_ram_111__1 (.Q (camera_module_cache_ram_111__1)
         , .QB (\$dummy [1301]), .D (nx3923), .CLK (clk), .R (rst)) ;
    mux21_ni ix3924 (.Y (nx3923), .A0 (nx35210), .A1 (
             camera_module_cache_ram_111__1), .S0 (nx36756)) ;
    nand04 ix6179 (.Y (nx6178), .A0 (nx29924), .A1 (nx29932), .A2 (nx29940), .A3 (
           nx29948)) ;
    aoi22 ix29925 (.Y (nx29924), .A0 (camera_module_cache_ram_143__1), .A1 (
          nx36150), .B0 (camera_module_cache_ram_159__1), .B1 (nx36190)) ;
    dffr camera_module_cache_reg_ram_143__1 (.Q (camera_module_cache_ram_143__1)
         , .QB (\$dummy [1302]), .D (nx3903), .CLK (clk), .R (rst)) ;
    mux21_ni ix3904 (.Y (nx3903), .A0 (nx35210), .A1 (
             camera_module_cache_ram_143__1), .S0 (nx36760)) ;
    dffr camera_module_cache_reg_ram_159__1 (.Q (camera_module_cache_ram_159__1)
         , .QB (\$dummy [1303]), .D (nx3893), .CLK (clk), .R (rst)) ;
    mux21_ni ix3894 (.Y (nx3893), .A0 (nx35210), .A1 (
             camera_module_cache_ram_159__1), .S0 (nx36764)) ;
    aoi22 ix29933 (.Y (nx29932), .A0 (camera_module_cache_ram_191__1), .A1 (
          nx36230), .B0 (camera_module_cache_ram_175__1), .B1 (nx36270)) ;
    dffr camera_module_cache_reg_ram_191__1 (.Q (camera_module_cache_ram_191__1)
         , .QB (\$dummy [1304]), .D (nx3873), .CLK (clk), .R (rst)) ;
    mux21_ni ix3874 (.Y (nx3873), .A0 (nx35210), .A1 (
             camera_module_cache_ram_191__1), .S0 (nx36768)) ;
    dffr camera_module_cache_reg_ram_175__1 (.Q (camera_module_cache_ram_175__1)
         , .QB (\$dummy [1305]), .D (nx3883), .CLK (clk), .R (rst)) ;
    mux21_ni ix3884 (.Y (nx3883), .A0 (nx35210), .A1 (
             camera_module_cache_ram_175__1), .S0 (nx36772)) ;
    aoi22 ix29941 (.Y (nx29940), .A0 (camera_module_cache_ram_207__1), .A1 (
          nx36310), .B0 (camera_module_cache_ram_223__1), .B1 (nx36350)) ;
    dffr camera_module_cache_reg_ram_207__1 (.Q (camera_module_cache_ram_207__1)
         , .QB (\$dummy [1306]), .D (nx3863), .CLK (clk), .R (rst)) ;
    mux21_ni ix3864 (.Y (nx3863), .A0 (nx35212), .A1 (
             camera_module_cache_ram_207__1), .S0 (nx36776)) ;
    dffr camera_module_cache_reg_ram_223__1 (.Q (camera_module_cache_ram_223__1)
         , .QB (\$dummy [1307]), .D (nx3853), .CLK (clk), .R (rst)) ;
    mux21_ni ix3854 (.Y (nx3853), .A0 (nx35212), .A1 (
             camera_module_cache_ram_223__1), .S0 (nx36780)) ;
    aoi22 ix29949 (.Y (nx29948), .A0 (camera_module_cache_ram_239__1), .A1 (
          nx36390), .B0 (camera_module_cache_ram_255__1), .B1 (nx36430)) ;
    dffr camera_module_cache_reg_ram_239__1 (.Q (camera_module_cache_ram_239__1)
         , .QB (\$dummy [1308]), .D (nx3843), .CLK (clk), .R (rst)) ;
    mux21_ni ix3844 (.Y (nx3843), .A0 (nx35212), .A1 (
             camera_module_cache_ram_239__1), .S0 (nx36784)) ;
    dffr camera_module_cache_reg_ram_255__1 (.Q (camera_module_cache_ram_255__1)
         , .QB (\$dummy [1309]), .D (nx3833), .CLK (clk), .R (rst)) ;
    mux21_ni ix3834 (.Y (nx3833), .A0 (nx35212), .A1 (
             camera_module_cache_ram_255__1), .S0 (nx36788)) ;
    dff camera_module_algo_module_pixel_reg_reg_q_3 (.Q (
        camera_module_algo_module_pixel_value_3), .QB (nx31098), .D (nx11533), .CLK (
        clk)) ;
    mux21_ni ix11534 (.Y (nx11533), .A0 (nx14286), .A1 (
             camera_module_algo_module_pixel_value_3), .S0 (nx22665)) ;
    mux21_ni ix29965 (.Y (nx29964), .A0 (nx29966), .A1 (nx35676), .S0 (nx36792)
             ) ;
    nor04 ix29967 (.Y (nx29966), .A0 (nx14266), .A1 (nx13612), .A2 (nx12956), .A3 (
          nx12302)) ;
    nand04 ix14267 (.Y (nx14266), .A0 (nx29969), .A1 (nx30075), .A2 (nx30143), .A3 (
           nx30211)) ;
    oai21 ix29970 (.Y (nx29969), .A0 (nx14256), .A1 (nx14178), .B0 (nx36448)) ;
    nand04 ix14257 (.Y (nx14256), .A0 (nx29972), .A1 (nx30018), .A2 (nx30026), .A3 (
           nx30034)) ;
    aoi22 ix29973 (.Y (nx29972), .A0 (camera_module_cache_ram_0__3), .A1 (
          nx35832), .B0 (camera_module_cache_ram_16__3), .B1 (nx35872)) ;
    dffr camera_module_cache_reg_ram_0__3 (.Q (camera_module_cache_ram_0__3), .QB (
         \$dummy [1310]), .D (nx11523), .CLK (clk), .R (rst)) ;
    mux21_ni ix11524 (.Y (nx11523), .A0 (camera_module_cache_ram_0__3), .A1 (
             nx35292), .S0 (nx35134)) ;
    oai221 ix11649 (.Y (nx11648), .A0 (nx34076), .A1 (nx29977), .B0 (nx29993), .B1 (
           nx35714), .C0 (nx29996)) ;
    tri01 nvm_module_tri_dataout_123 (.Y (nvm_data_123), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_115 (.Y (nvm_data_115), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_107 (.Y (nvm_data_107), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_99 (.Y (nvm_data_99), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_91 (.Y (nvm_data_91), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_83 (.Y (nvm_data_83), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_75 (.Y (nvm_data_75), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_67 (.Y (nvm_data_67), .A (nx22549), .E (
          nvm_module_GND0)) ;
    inv01 ix29994 (.Y (nx29993), .A (nvm_data_3)) ;
    tri01 nvm_module_tri_dataout_3 (.Y (nvm_data_3), .A (nx22549), .E (
          nvm_module_GND0)) ;
    nand02 ix29997 (.Y (nx29996), .A0 (nx34076), .A1 (nx11582)) ;
    tri01 nvm_module_tri_dataout_59 (.Y (nvm_data_59), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_51 (.Y (nvm_data_51), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_43 (.Y (nvm_data_43), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_35 (.Y (nvm_data_35), .A (nx22549), .E (
          nvm_module_GND0)) ;
    oai22 ix11551 (.Y (nx11550), .A0 (nx34106), .A1 (nx30007), .B0 (nx34092), .B1 (
          nx30011)) ;
    tri01 nvm_module_tri_dataout_27 (.Y (nvm_data_27), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_19 (.Y (nvm_data_19), .A (nx22549), .E (
          nvm_module_GND0)) ;
    nand02 ix30012 (.Y (nx30011), .A0 (nvm_data_11), .A1 (nx34106)) ;
    tri01 nvm_module_tri_dataout_11 (.Y (nvm_data_11), .A (nx22549), .E (
          nvm_module_GND0)) ;
    dffr camera_module_cache_reg_ram_16__3 (.Q (camera_module_cache_ram_16__3), 
         .QB (\$dummy [1311]), .D (nx11513), .CLK (clk), .R (rst)) ;
    mux21_ni ix11514 (.Y (nx11513), .A0 (camera_module_cache_ram_16__3), .A1 (
             nx35292), .S0 (nx35130)) ;
    aoi22 ix30019 (.Y (nx30018), .A0 (camera_module_cache_ram_32__3), .A1 (
          nx35912), .B0 (camera_module_cache_ram_48__3), .B1 (nx35952)) ;
    dffr camera_module_cache_reg_ram_32__3 (.Q (camera_module_cache_ram_32__3), 
         .QB (\$dummy [1312]), .D (nx11503), .CLK (clk), .R (rst)) ;
    mux21_ni ix11504 (.Y (nx11503), .A0 (camera_module_cache_ram_32__3), .A1 (
             nx35292), .S0 (nx35126)) ;
    dffr camera_module_cache_reg_ram_48__3 (.Q (camera_module_cache_ram_48__3), 
         .QB (\$dummy [1313]), .D (nx11493), .CLK (clk), .R (rst)) ;
    mux21_ni ix11494 (.Y (nx11493), .A0 (camera_module_cache_ram_48__3), .A1 (
             nx35292), .S0 (nx35122)) ;
    aoi22 ix30027 (.Y (nx30026), .A0 (camera_module_cache_ram_64__3), .A1 (
          nx35992), .B0 (camera_module_cache_ram_80__3), .B1 (nx36032)) ;
    dffr camera_module_cache_reg_ram_64__3 (.Q (camera_module_cache_ram_64__3), 
         .QB (\$dummy [1314]), .D (nx11483), .CLK (clk), .R (rst)) ;
    mux21_ni ix11484 (.Y (nx11483), .A0 (camera_module_cache_ram_64__3), .A1 (
             nx35292), .S0 (nx35118)) ;
    dffr camera_module_cache_reg_ram_80__3 (.Q (camera_module_cache_ram_80__3), 
         .QB (\$dummy [1315]), .D (nx11473), .CLK (clk), .R (rst)) ;
    mux21_ni ix11474 (.Y (nx11473), .A0 (camera_module_cache_ram_80__3), .A1 (
             nx35292), .S0 (nx35114)) ;
    aoi22 ix30035 (.Y (nx30034), .A0 (camera_module_cache_ram_112__3), .A1 (
          nx36072), .B0 (camera_module_cache_ram_96__3), .B1 (nx36112)) ;
    dffr camera_module_cache_reg_ram_112__3 (.Q (camera_module_cache_ram_112__3)
         , .QB (\$dummy [1316]), .D (nx11453), .CLK (clk), .R (rst)) ;
    mux21_ni ix11454 (.Y (nx11453), .A0 (camera_module_cache_ram_112__3), .A1 (
             nx35292), .S0 (nx35106)) ;
    dffr camera_module_cache_reg_ram_96__3 (.Q (camera_module_cache_ram_96__3), 
         .QB (\$dummy [1317]), .D (nx11463), .CLK (clk), .R (rst)) ;
    mux21_ni ix11464 (.Y (nx11463), .A0 (camera_module_cache_ram_96__3), .A1 (
             nx35294), .S0 (nx35110)) ;
    nand04 ix14179 (.Y (nx14178), .A0 (nx30043), .A1 (nx30051), .A2 (nx30059), .A3 (
           nx30067)) ;
    aoi22 ix30044 (.Y (nx30043), .A0 (camera_module_cache_ram_128__3), .A1 (
          nx36152), .B0 (camera_module_cache_ram_144__3), .B1 (nx36192)) ;
    dffr camera_module_cache_reg_ram_128__3 (.Q (camera_module_cache_ram_128__3)
         , .QB (\$dummy [1318]), .D (nx11443), .CLK (clk), .R (rst)) ;
    mux21_ni ix11444 (.Y (nx11443), .A0 (camera_module_cache_ram_128__3), .A1 (
             nx35294), .S0 (nx35102)) ;
    dffr camera_module_cache_reg_ram_144__3 (.Q (camera_module_cache_ram_144__3)
         , .QB (\$dummy [1319]), .D (nx11433), .CLK (clk), .R (rst)) ;
    mux21_ni ix11434 (.Y (nx11433), .A0 (camera_module_cache_ram_144__3), .A1 (
             nx35294), .S0 (nx35098)) ;
    aoi22 ix30052 (.Y (nx30051), .A0 (camera_module_cache_ram_176__3), .A1 (
          nx36232), .B0 (camera_module_cache_ram_160__3), .B1 (nx36272)) ;
    dffr camera_module_cache_reg_ram_176__3 (.Q (camera_module_cache_ram_176__3)
         , .QB (\$dummy [1320]), .D (nx11413), .CLK (clk), .R (rst)) ;
    mux21_ni ix11414 (.Y (nx11413), .A0 (camera_module_cache_ram_176__3), .A1 (
             nx35294), .S0 (nx35090)) ;
    dffr camera_module_cache_reg_ram_160__3 (.Q (camera_module_cache_ram_160__3)
         , .QB (\$dummy [1321]), .D (nx11423), .CLK (clk), .R (rst)) ;
    mux21_ni ix11424 (.Y (nx11423), .A0 (camera_module_cache_ram_160__3), .A1 (
             nx35294), .S0 (nx35094)) ;
    aoi22 ix30060 (.Y (nx30059), .A0 (camera_module_cache_ram_192__3), .A1 (
          nx36312), .B0 (camera_module_cache_ram_208__3), .B1 (nx36352)) ;
    dffr camera_module_cache_reg_ram_192__3 (.Q (camera_module_cache_ram_192__3)
         , .QB (\$dummy [1322]), .D (nx11403), .CLK (clk), .R (rst)) ;
    mux21_ni ix11404 (.Y (nx11403), .A0 (camera_module_cache_ram_192__3), .A1 (
             nx35294), .S0 (nx35086)) ;
    dffr camera_module_cache_reg_ram_208__3 (.Q (camera_module_cache_ram_208__3)
         , .QB (\$dummy [1323]), .D (nx11393), .CLK (clk), .R (rst)) ;
    mux21_ni ix11394 (.Y (nx11393), .A0 (camera_module_cache_ram_208__3), .A1 (
             nx35294), .S0 (nx35082)) ;
    aoi22 ix30068 (.Y (nx30067), .A0 (camera_module_cache_ram_224__3), .A1 (
          nx36392), .B0 (camera_module_cache_ram_240__3), .B1 (nx36432)) ;
    dffr camera_module_cache_reg_ram_224__3 (.Q (camera_module_cache_ram_224__3)
         , .QB (\$dummy [1324]), .D (nx11383), .CLK (clk), .R (rst)) ;
    mux21_ni ix11384 (.Y (nx11383), .A0 (camera_module_cache_ram_224__3), .A1 (
             nx35296), .S0 (nx35078)) ;
    dffr camera_module_cache_reg_ram_240__3 (.Q (camera_module_cache_ram_240__3)
         , .QB (\$dummy [1325]), .D (nx11373), .CLK (clk), .R (rst)) ;
    mux21_ni ix11374 (.Y (nx11373), .A0 (camera_module_cache_ram_240__3), .A1 (
             nx35296), .S0 (nx35074)) ;
    oai21 ix30076 (.Y (nx30075), .A0 (nx14094), .A1 (nx14016), .B0 (nx36452)) ;
    nand04 ix14095 (.Y (nx14094), .A0 (nx30078), .A1 (nx30086), .A2 (nx30094), .A3 (
           nx30102)) ;
    aoi22 ix30079 (.Y (nx30078), .A0 (camera_module_cache_ram_1__3), .A1 (
          nx35832), .B0 (camera_module_cache_ram_17__3), .B1 (nx35872)) ;
    dffr camera_module_cache_reg_ram_1__3 (.Q (camera_module_cache_ram_1__3), .QB (
         \$dummy [1326]), .D (nx11363), .CLK (clk), .R (rst)) ;
    mux21_ni ix11364 (.Y (nx11363), .A0 (camera_module_cache_ram_1__3), .A1 (
             nx35296), .S0 (nx35064)) ;
    dffr camera_module_cache_reg_ram_17__3 (.Q (camera_module_cache_ram_17__3), 
         .QB (\$dummy [1327]), .D (nx11353), .CLK (clk), .R (rst)) ;
    mux21_ni ix11354 (.Y (nx11353), .A0 (camera_module_cache_ram_17__3), .A1 (
             nx35296), .S0 (nx35060)) ;
    aoi22 ix30087 (.Y (nx30086), .A0 (camera_module_cache_ram_33__3), .A1 (
          nx35912), .B0 (camera_module_cache_ram_49__3), .B1 (nx35952)) ;
    dffr camera_module_cache_reg_ram_33__3 (.Q (camera_module_cache_ram_33__3), 
         .QB (\$dummy [1328]), .D (nx11343), .CLK (clk), .R (rst)) ;
    mux21_ni ix11344 (.Y (nx11343), .A0 (camera_module_cache_ram_33__3), .A1 (
             nx35296), .S0 (nx35056)) ;
    dffr camera_module_cache_reg_ram_49__3 (.Q (camera_module_cache_ram_49__3), 
         .QB (\$dummy [1329]), .D (nx11333), .CLK (clk), .R (rst)) ;
    mux21_ni ix11334 (.Y (nx11333), .A0 (camera_module_cache_ram_49__3), .A1 (
             nx35296), .S0 (nx35052)) ;
    aoi22 ix30095 (.Y (nx30094), .A0 (camera_module_cache_ram_65__3), .A1 (
          nx35992), .B0 (camera_module_cache_ram_81__3), .B1 (nx36032)) ;
    dffr camera_module_cache_reg_ram_65__3 (.Q (camera_module_cache_ram_65__3), 
         .QB (\$dummy [1330]), .D (nx11323), .CLK (clk), .R (rst)) ;
    mux21_ni ix11324 (.Y (nx11323), .A0 (camera_module_cache_ram_65__3), .A1 (
             nx35296), .S0 (nx35048)) ;
    dffr camera_module_cache_reg_ram_81__3 (.Q (camera_module_cache_ram_81__3), 
         .QB (\$dummy [1331]), .D (nx11313), .CLK (clk), .R (rst)) ;
    mux21_ni ix11314 (.Y (nx11313), .A0 (camera_module_cache_ram_81__3), .A1 (
             nx35298), .S0 (nx35044)) ;
    aoi22 ix30103 (.Y (nx30102), .A0 (camera_module_cache_ram_113__3), .A1 (
          nx36072), .B0 (camera_module_cache_ram_97__3), .B1 (nx36112)) ;
    dffr camera_module_cache_reg_ram_113__3 (.Q (camera_module_cache_ram_113__3)
         , .QB (\$dummy [1332]), .D (nx11293), .CLK (clk), .R (rst)) ;
    mux21_ni ix11294 (.Y (nx11293), .A0 (camera_module_cache_ram_113__3), .A1 (
             nx35298), .S0 (nx35036)) ;
    dffr camera_module_cache_reg_ram_97__3 (.Q (camera_module_cache_ram_97__3), 
         .QB (\$dummy [1333]), .D (nx11303), .CLK (clk), .R (rst)) ;
    mux21_ni ix11304 (.Y (nx11303), .A0 (camera_module_cache_ram_97__3), .A1 (
             nx35298), .S0 (nx35040)) ;
    nand04 ix14017 (.Y (nx14016), .A0 (nx30111), .A1 (nx30119), .A2 (nx30127), .A3 (
           nx30135)) ;
    aoi22 ix30112 (.Y (nx30111), .A0 (camera_module_cache_ram_129__3), .A1 (
          nx36152), .B0 (camera_module_cache_ram_145__3), .B1 (nx36192)) ;
    dffr camera_module_cache_reg_ram_129__3 (.Q (camera_module_cache_ram_129__3)
         , .QB (\$dummy [1334]), .D (nx11283), .CLK (clk), .R (rst)) ;
    mux21_ni ix11284 (.Y (nx11283), .A0 (camera_module_cache_ram_129__3), .A1 (
             nx35298), .S0 (nx35032)) ;
    dffr camera_module_cache_reg_ram_145__3 (.Q (camera_module_cache_ram_145__3)
         , .QB (\$dummy [1335]), .D (nx11273), .CLK (clk), .R (rst)) ;
    mux21_ni ix11274 (.Y (nx11273), .A0 (camera_module_cache_ram_145__3), .A1 (
             nx35298), .S0 (nx35028)) ;
    aoi22 ix30120 (.Y (nx30119), .A0 (camera_module_cache_ram_177__3), .A1 (
          nx36232), .B0 (camera_module_cache_ram_161__3), .B1 (nx36272)) ;
    dffr camera_module_cache_reg_ram_177__3 (.Q (camera_module_cache_ram_177__3)
         , .QB (\$dummy [1336]), .D (nx11253), .CLK (clk), .R (rst)) ;
    mux21_ni ix11254 (.Y (nx11253), .A0 (camera_module_cache_ram_177__3), .A1 (
             nx35298), .S0 (nx35020)) ;
    dffr camera_module_cache_reg_ram_161__3 (.Q (camera_module_cache_ram_161__3)
         , .QB (\$dummy [1337]), .D (nx11263), .CLK (clk), .R (rst)) ;
    mux21_ni ix11264 (.Y (nx11263), .A0 (camera_module_cache_ram_161__3), .A1 (
             nx35298), .S0 (nx35024)) ;
    aoi22 ix30128 (.Y (nx30127), .A0 (camera_module_cache_ram_193__3), .A1 (
          nx36312), .B0 (camera_module_cache_ram_209__3), .B1 (nx36352)) ;
    dffr camera_module_cache_reg_ram_193__3 (.Q (camera_module_cache_ram_193__3)
         , .QB (\$dummy [1338]), .D (nx11243), .CLK (clk), .R (rst)) ;
    mux21_ni ix11244 (.Y (nx11243), .A0 (camera_module_cache_ram_193__3), .A1 (
             nx35300), .S0 (nx35016)) ;
    dffr camera_module_cache_reg_ram_209__3 (.Q (camera_module_cache_ram_209__3)
         , .QB (\$dummy [1339]), .D (nx11233), .CLK (clk), .R (rst)) ;
    mux21_ni ix11234 (.Y (nx11233), .A0 (camera_module_cache_ram_209__3), .A1 (
             nx35300), .S0 (nx35012)) ;
    aoi22 ix30136 (.Y (nx30135), .A0 (camera_module_cache_ram_225__3), .A1 (
          nx36392), .B0 (camera_module_cache_ram_241__3), .B1 (nx36432)) ;
    dffr camera_module_cache_reg_ram_225__3 (.Q (camera_module_cache_ram_225__3)
         , .QB (\$dummy [1340]), .D (nx11223), .CLK (clk), .R (rst)) ;
    mux21_ni ix11224 (.Y (nx11223), .A0 (camera_module_cache_ram_225__3), .A1 (
             nx35300), .S0 (nx35008)) ;
    dffr camera_module_cache_reg_ram_241__3 (.Q (camera_module_cache_ram_241__3)
         , .QB (\$dummy [1341]), .D (nx11213), .CLK (clk), .R (rst)) ;
    mux21_ni ix11214 (.Y (nx11213), .A0 (camera_module_cache_ram_241__3), .A1 (
             nx35300), .S0 (nx35004)) ;
    oai21 ix30144 (.Y (nx30143), .A0 (nx13930), .A1 (nx13852), .B0 (nx36456)) ;
    nand04 ix13931 (.Y (nx13930), .A0 (nx30146), .A1 (nx30154), .A2 (nx30162), .A3 (
           nx30170)) ;
    aoi22 ix30147 (.Y (nx30146), .A0 (camera_module_cache_ram_2__3), .A1 (
          nx35832), .B0 (camera_module_cache_ram_18__3), .B1 (nx35872)) ;
    dffr camera_module_cache_reg_ram_2__3 (.Q (camera_module_cache_ram_2__3), .QB (
         \$dummy [1342]), .D (nx11203), .CLK (clk), .R (rst)) ;
    mux21_ni ix11204 (.Y (nx11203), .A0 (camera_module_cache_ram_2__3), .A1 (
             nx35300), .S0 (nx34994)) ;
    dffr camera_module_cache_reg_ram_18__3 (.Q (camera_module_cache_ram_18__3), 
         .QB (\$dummy [1343]), .D (nx11193), .CLK (clk), .R (rst)) ;
    mux21_ni ix11194 (.Y (nx11193), .A0 (camera_module_cache_ram_18__3), .A1 (
             nx35300), .S0 (nx34990)) ;
    aoi22 ix30155 (.Y (nx30154), .A0 (camera_module_cache_ram_34__3), .A1 (
          nx35912), .B0 (camera_module_cache_ram_50__3), .B1 (nx35952)) ;
    dffr camera_module_cache_reg_ram_34__3 (.Q (camera_module_cache_ram_34__3), 
         .QB (\$dummy [1344]), .D (nx11183), .CLK (clk), .R (rst)) ;
    mux21_ni ix11184 (.Y (nx11183), .A0 (camera_module_cache_ram_34__3), .A1 (
             nx35300), .S0 (nx34986)) ;
    dffr camera_module_cache_reg_ram_50__3 (.Q (camera_module_cache_ram_50__3), 
         .QB (\$dummy [1345]), .D (nx11173), .CLK (clk), .R (rst)) ;
    mux21_ni ix11174 (.Y (nx11173), .A0 (camera_module_cache_ram_50__3), .A1 (
             nx35302), .S0 (nx34982)) ;
    aoi22 ix30163 (.Y (nx30162), .A0 (camera_module_cache_ram_66__3), .A1 (
          nx35992), .B0 (camera_module_cache_ram_82__3), .B1 (nx36032)) ;
    dffr camera_module_cache_reg_ram_66__3 (.Q (camera_module_cache_ram_66__3), 
         .QB (\$dummy [1346]), .D (nx11163), .CLK (clk), .R (rst)) ;
    mux21_ni ix11164 (.Y (nx11163), .A0 (camera_module_cache_ram_66__3), .A1 (
             nx35302), .S0 (nx34978)) ;
    dffr camera_module_cache_reg_ram_82__3 (.Q (camera_module_cache_ram_82__3), 
         .QB (\$dummy [1347]), .D (nx11153), .CLK (clk), .R (rst)) ;
    mux21_ni ix11154 (.Y (nx11153), .A0 (camera_module_cache_ram_82__3), .A1 (
             nx35302), .S0 (nx34974)) ;
    aoi22 ix30171 (.Y (nx30170), .A0 (camera_module_cache_ram_114__3), .A1 (
          nx36072), .B0 (camera_module_cache_ram_98__3), .B1 (nx36112)) ;
    dffr camera_module_cache_reg_ram_114__3 (.Q (camera_module_cache_ram_114__3)
         , .QB (\$dummy [1348]), .D (nx11133), .CLK (clk), .R (rst)) ;
    mux21_ni ix11134 (.Y (nx11133), .A0 (camera_module_cache_ram_114__3), .A1 (
             nx35302), .S0 (nx34966)) ;
    dffr camera_module_cache_reg_ram_98__3 (.Q (camera_module_cache_ram_98__3), 
         .QB (\$dummy [1349]), .D (nx11143), .CLK (clk), .R (rst)) ;
    mux21_ni ix11144 (.Y (nx11143), .A0 (camera_module_cache_ram_98__3), .A1 (
             nx35302), .S0 (nx34970)) ;
    nand04 ix13853 (.Y (nx13852), .A0 (nx30179), .A1 (nx30187), .A2 (nx30195), .A3 (
           nx30203)) ;
    aoi22 ix30180 (.Y (nx30179), .A0 (camera_module_cache_ram_130__3), .A1 (
          nx36152), .B0 (camera_module_cache_ram_146__3), .B1 (nx36192)) ;
    dffr camera_module_cache_reg_ram_130__3 (.Q (camera_module_cache_ram_130__3)
         , .QB (\$dummy [1350]), .D (nx11123), .CLK (clk), .R (rst)) ;
    mux21_ni ix11124 (.Y (nx11123), .A0 (camera_module_cache_ram_130__3), .A1 (
             nx35302), .S0 (nx34962)) ;
    dffr camera_module_cache_reg_ram_146__3 (.Q (camera_module_cache_ram_146__3)
         , .QB (\$dummy [1351]), .D (nx11113), .CLK (clk), .R (rst)) ;
    mux21_ni ix11114 (.Y (nx11113), .A0 (camera_module_cache_ram_146__3), .A1 (
             nx35302), .S0 (nx34958)) ;
    aoi22 ix30188 (.Y (nx30187), .A0 (camera_module_cache_ram_178__3), .A1 (
          nx36232), .B0 (camera_module_cache_ram_162__3), .B1 (nx36272)) ;
    dffr camera_module_cache_reg_ram_178__3 (.Q (camera_module_cache_ram_178__3)
         , .QB (\$dummy [1352]), .D (nx11093), .CLK (clk), .R (rst)) ;
    mux21_ni ix11094 (.Y (nx11093), .A0 (camera_module_cache_ram_178__3), .A1 (
             nx35304), .S0 (nx34950)) ;
    dffr camera_module_cache_reg_ram_162__3 (.Q (camera_module_cache_ram_162__3)
         , .QB (\$dummy [1353]), .D (nx11103), .CLK (clk), .R (rst)) ;
    mux21_ni ix11104 (.Y (nx11103), .A0 (camera_module_cache_ram_162__3), .A1 (
             nx35304), .S0 (nx34954)) ;
    aoi22 ix30196 (.Y (nx30195), .A0 (camera_module_cache_ram_194__3), .A1 (
          nx36312), .B0 (camera_module_cache_ram_210__3), .B1 (nx36352)) ;
    dffr camera_module_cache_reg_ram_194__3 (.Q (camera_module_cache_ram_194__3)
         , .QB (\$dummy [1354]), .D (nx11083), .CLK (clk), .R (rst)) ;
    mux21_ni ix11084 (.Y (nx11083), .A0 (camera_module_cache_ram_194__3), .A1 (
             nx35304), .S0 (nx34946)) ;
    dffr camera_module_cache_reg_ram_210__3 (.Q (camera_module_cache_ram_210__3)
         , .QB (\$dummy [1355]), .D (nx11073), .CLK (clk), .R (rst)) ;
    mux21_ni ix11074 (.Y (nx11073), .A0 (camera_module_cache_ram_210__3), .A1 (
             nx35304), .S0 (nx34942)) ;
    aoi22 ix30204 (.Y (nx30203), .A0 (camera_module_cache_ram_226__3), .A1 (
          nx36392), .B0 (camera_module_cache_ram_242__3), .B1 (nx36432)) ;
    dffr camera_module_cache_reg_ram_226__3 (.Q (camera_module_cache_ram_226__3)
         , .QB (\$dummy [1356]), .D (nx11063), .CLK (clk), .R (rst)) ;
    mux21_ni ix11064 (.Y (nx11063), .A0 (camera_module_cache_ram_226__3), .A1 (
             nx35304), .S0 (nx34938)) ;
    dffr camera_module_cache_reg_ram_242__3 (.Q (camera_module_cache_ram_242__3)
         , .QB (\$dummy [1357]), .D (nx11053), .CLK (clk), .R (rst)) ;
    mux21_ni ix11054 (.Y (nx11053), .A0 (camera_module_cache_ram_242__3), .A1 (
             nx35304), .S0 (nx34934)) ;
    oai21 ix30212 (.Y (nx30211), .A0 (nx13768), .A1 (nx13690), .B0 (nx36460)) ;
    nand04 ix13769 (.Y (nx13768), .A0 (nx30214), .A1 (nx30222), .A2 (nx30230), .A3 (
           nx30238)) ;
    aoi22 ix30215 (.Y (nx30214), .A0 (camera_module_cache_ram_3__3), .A1 (
          nx35832), .B0 (camera_module_cache_ram_19__3), .B1 (nx35872)) ;
    dffr camera_module_cache_reg_ram_3__3 (.Q (camera_module_cache_ram_3__3), .QB (
         \$dummy [1358]), .D (nx11043), .CLK (clk), .R (rst)) ;
    mux21_ni ix11044 (.Y (nx11043), .A0 (camera_module_cache_ram_3__3), .A1 (
             nx35304), .S0 (nx34924)) ;
    dffr camera_module_cache_reg_ram_19__3 (.Q (camera_module_cache_ram_19__3), 
         .QB (\$dummy [1359]), .D (nx11033), .CLK (clk), .R (rst)) ;
    mux21_ni ix11034 (.Y (nx11033), .A0 (camera_module_cache_ram_19__3), .A1 (
             nx35306), .S0 (nx34920)) ;
    aoi22 ix30223 (.Y (nx30222), .A0 (camera_module_cache_ram_35__3), .A1 (
          nx35912), .B0 (camera_module_cache_ram_51__3), .B1 (nx35952)) ;
    dffr camera_module_cache_reg_ram_35__3 (.Q (camera_module_cache_ram_35__3), 
         .QB (\$dummy [1360]), .D (nx11023), .CLK (clk), .R (rst)) ;
    mux21_ni ix11024 (.Y (nx11023), .A0 (camera_module_cache_ram_35__3), .A1 (
             nx35306), .S0 (nx34916)) ;
    dffr camera_module_cache_reg_ram_51__3 (.Q (camera_module_cache_ram_51__3), 
         .QB (\$dummy [1361]), .D (nx11013), .CLK (clk), .R (rst)) ;
    mux21_ni ix11014 (.Y (nx11013), .A0 (camera_module_cache_ram_51__3), .A1 (
             nx35306), .S0 (nx34912)) ;
    aoi22 ix30231 (.Y (nx30230), .A0 (camera_module_cache_ram_67__3), .A1 (
          nx35992), .B0 (camera_module_cache_ram_83__3), .B1 (nx36032)) ;
    dffr camera_module_cache_reg_ram_67__3 (.Q (camera_module_cache_ram_67__3), 
         .QB (\$dummy [1362]), .D (nx11003), .CLK (clk), .R (rst)) ;
    mux21_ni ix11004 (.Y (nx11003), .A0 (camera_module_cache_ram_67__3), .A1 (
             nx35306), .S0 (nx34908)) ;
    dffr camera_module_cache_reg_ram_83__3 (.Q (camera_module_cache_ram_83__3), 
         .QB (\$dummy [1363]), .D (nx10993), .CLK (clk), .R (rst)) ;
    mux21_ni ix10994 (.Y (nx10993), .A0 (camera_module_cache_ram_83__3), .A1 (
             nx35306), .S0 (nx34904)) ;
    aoi22 ix30239 (.Y (nx30238), .A0 (camera_module_cache_ram_115__3), .A1 (
          nx36072), .B0 (camera_module_cache_ram_99__3), .B1 (nx36112)) ;
    dffr camera_module_cache_reg_ram_115__3 (.Q (camera_module_cache_ram_115__3)
         , .QB (\$dummy [1364]), .D (nx10973), .CLK (clk), .R (rst)) ;
    mux21_ni ix10974 (.Y (nx10973), .A0 (camera_module_cache_ram_115__3), .A1 (
             nx35306), .S0 (nx34896)) ;
    dffr camera_module_cache_reg_ram_99__3 (.Q (camera_module_cache_ram_99__3), 
         .QB (\$dummy [1365]), .D (nx10983), .CLK (clk), .R (rst)) ;
    mux21_ni ix10984 (.Y (nx10983), .A0 (camera_module_cache_ram_99__3), .A1 (
             nx35306), .S0 (nx34900)) ;
    nand04 ix13691 (.Y (nx13690), .A0 (nx30247), .A1 (nx30255), .A2 (nx30263), .A3 (
           nx30271)) ;
    aoi22 ix30248 (.Y (nx30247), .A0 (camera_module_cache_ram_131__3), .A1 (
          nx36152), .B0 (camera_module_cache_ram_147__3), .B1 (nx36192)) ;
    dffr camera_module_cache_reg_ram_131__3 (.Q (camera_module_cache_ram_131__3)
         , .QB (\$dummy [1366]), .D (nx10963), .CLK (clk), .R (rst)) ;
    mux21_ni ix10964 (.Y (nx10963), .A0 (camera_module_cache_ram_131__3), .A1 (
             nx35308), .S0 (nx34892)) ;
    dffr camera_module_cache_reg_ram_147__3 (.Q (camera_module_cache_ram_147__3)
         , .QB (\$dummy [1367]), .D (nx10953), .CLK (clk), .R (rst)) ;
    mux21_ni ix10954 (.Y (nx10953), .A0 (camera_module_cache_ram_147__3), .A1 (
             nx35308), .S0 (nx34888)) ;
    aoi22 ix30256 (.Y (nx30255), .A0 (camera_module_cache_ram_179__3), .A1 (
          nx36232), .B0 (camera_module_cache_ram_163__3), .B1 (nx36272)) ;
    dffr camera_module_cache_reg_ram_179__3 (.Q (camera_module_cache_ram_179__3)
         , .QB (\$dummy [1368]), .D (nx10933), .CLK (clk), .R (rst)) ;
    mux21_ni ix10934 (.Y (nx10933), .A0 (camera_module_cache_ram_179__3), .A1 (
             nx35308), .S0 (nx34880)) ;
    dffr camera_module_cache_reg_ram_163__3 (.Q (camera_module_cache_ram_163__3)
         , .QB (\$dummy [1369]), .D (nx10943), .CLK (clk), .R (rst)) ;
    mux21_ni ix10944 (.Y (nx10943), .A0 (camera_module_cache_ram_163__3), .A1 (
             nx35308), .S0 (nx34884)) ;
    aoi22 ix30264 (.Y (nx30263), .A0 (camera_module_cache_ram_195__3), .A1 (
          nx36312), .B0 (camera_module_cache_ram_211__3), .B1 (nx36352)) ;
    dffr camera_module_cache_reg_ram_195__3 (.Q (camera_module_cache_ram_195__3)
         , .QB (\$dummy [1370]), .D (nx10923), .CLK (clk), .R (rst)) ;
    mux21_ni ix10924 (.Y (nx10923), .A0 (camera_module_cache_ram_195__3), .A1 (
             nx35308), .S0 (nx34876)) ;
    dffr camera_module_cache_reg_ram_211__3 (.Q (camera_module_cache_ram_211__3)
         , .QB (\$dummy [1371]), .D (nx10913), .CLK (clk), .R (rst)) ;
    mux21_ni ix10914 (.Y (nx10913), .A0 (camera_module_cache_ram_211__3), .A1 (
             nx35308), .S0 (nx34872)) ;
    aoi22 ix30272 (.Y (nx30271), .A0 (camera_module_cache_ram_227__3), .A1 (
          nx36392), .B0 (camera_module_cache_ram_243__3), .B1 (nx36432)) ;
    dffr camera_module_cache_reg_ram_227__3 (.Q (camera_module_cache_ram_227__3)
         , .QB (\$dummy [1372]), .D (nx10903), .CLK (clk), .R (rst)) ;
    mux21_ni ix10904 (.Y (nx10903), .A0 (camera_module_cache_ram_227__3), .A1 (
             nx35308), .S0 (nx34868)) ;
    dffr camera_module_cache_reg_ram_243__3 (.Q (camera_module_cache_ram_243__3)
         , .QB (\$dummy [1373]), .D (nx10893), .CLK (clk), .R (rst)) ;
    mux21_ni ix10894 (.Y (nx10893), .A0 (camera_module_cache_ram_243__3), .A1 (
             nx35310), .S0 (nx34864)) ;
    nand04 ix13613 (.Y (nx13612), .A0 (nx30280), .A1 (nx30348), .A2 (nx30416), .A3 (
           nx30484)) ;
    oai21 ix30281 (.Y (nx30280), .A0 (nx13602), .A1 (nx13524), .B0 (nx36464)) ;
    nand04 ix13603 (.Y (nx13602), .A0 (nx30283), .A1 (nx30291), .A2 (nx30299), .A3 (
           nx30307)) ;
    aoi22 ix30284 (.Y (nx30283), .A0 (camera_module_cache_ram_4__3), .A1 (
          nx35832), .B0 (camera_module_cache_ram_20__3), .B1 (nx35872)) ;
    dffr camera_module_cache_reg_ram_4__3 (.Q (camera_module_cache_ram_4__3), .QB (
         \$dummy [1374]), .D (nx10883), .CLK (clk), .R (rst)) ;
    mux21_ni ix10884 (.Y (nx10883), .A0 (camera_module_cache_ram_4__3), .A1 (
             nx35310), .S0 (nx34854)) ;
    dffr camera_module_cache_reg_ram_20__3 (.Q (camera_module_cache_ram_20__3), 
         .QB (\$dummy [1375]), .D (nx10873), .CLK (clk), .R (rst)) ;
    mux21_ni ix10874 (.Y (nx10873), .A0 (camera_module_cache_ram_20__3), .A1 (
             nx35310), .S0 (nx34850)) ;
    aoi22 ix30292 (.Y (nx30291), .A0 (camera_module_cache_ram_36__3), .A1 (
          nx35912), .B0 (camera_module_cache_ram_52__3), .B1 (nx35952)) ;
    dffr camera_module_cache_reg_ram_36__3 (.Q (camera_module_cache_ram_36__3), 
         .QB (\$dummy [1376]), .D (nx10863), .CLK (clk), .R (rst)) ;
    mux21_ni ix10864 (.Y (nx10863), .A0 (camera_module_cache_ram_36__3), .A1 (
             nx35310), .S0 (nx34846)) ;
    dffr camera_module_cache_reg_ram_52__3 (.Q (camera_module_cache_ram_52__3), 
         .QB (\$dummy [1377]), .D (nx10853), .CLK (clk), .R (rst)) ;
    mux21_ni ix10854 (.Y (nx10853), .A0 (camera_module_cache_ram_52__3), .A1 (
             nx35310), .S0 (nx34842)) ;
    aoi22 ix30300 (.Y (nx30299), .A0 (camera_module_cache_ram_68__3), .A1 (
          nx35992), .B0 (camera_module_cache_ram_84__3), .B1 (nx36032)) ;
    dffr camera_module_cache_reg_ram_68__3 (.Q (camera_module_cache_ram_68__3), 
         .QB (\$dummy [1378]), .D (nx10843), .CLK (clk), .R (rst)) ;
    mux21_ni ix10844 (.Y (nx10843), .A0 (camera_module_cache_ram_68__3), .A1 (
             nx35310), .S0 (nx34838)) ;
    dffr camera_module_cache_reg_ram_84__3 (.Q (camera_module_cache_ram_84__3), 
         .QB (\$dummy [1379]), .D (nx10833), .CLK (clk), .R (rst)) ;
    mux21_ni ix10834 (.Y (nx10833), .A0 (camera_module_cache_ram_84__3), .A1 (
             nx35310), .S0 (nx34834)) ;
    aoi22 ix30308 (.Y (nx30307), .A0 (camera_module_cache_ram_116__3), .A1 (
          nx36072), .B0 (camera_module_cache_ram_100__3), .B1 (nx36112)) ;
    dffr camera_module_cache_reg_ram_116__3 (.Q (camera_module_cache_ram_116__3)
         , .QB (\$dummy [1380]), .D (nx10813), .CLK (clk), .R (rst)) ;
    mux21_ni ix10814 (.Y (nx10813), .A0 (camera_module_cache_ram_116__3), .A1 (
             nx35312), .S0 (nx34826)) ;
    dffr camera_module_cache_reg_ram_100__3 (.Q (camera_module_cache_ram_100__3)
         , .QB (\$dummy [1381]), .D (nx10823), .CLK (clk), .R (rst)) ;
    mux21_ni ix10824 (.Y (nx10823), .A0 (camera_module_cache_ram_100__3), .A1 (
             nx35312), .S0 (nx34830)) ;
    nand04 ix13525 (.Y (nx13524), .A0 (nx30316), .A1 (nx30324), .A2 (nx30332), .A3 (
           nx30340)) ;
    aoi22 ix30317 (.Y (nx30316), .A0 (camera_module_cache_ram_132__3), .A1 (
          nx36152), .B0 (camera_module_cache_ram_148__3), .B1 (nx36192)) ;
    dffr camera_module_cache_reg_ram_132__3 (.Q (camera_module_cache_ram_132__3)
         , .QB (\$dummy [1382]), .D (nx10803), .CLK (clk), .R (rst)) ;
    mux21_ni ix10804 (.Y (nx10803), .A0 (camera_module_cache_ram_132__3), .A1 (
             nx35312), .S0 (nx34822)) ;
    dffr camera_module_cache_reg_ram_148__3 (.Q (camera_module_cache_ram_148__3)
         , .QB (\$dummy [1383]), .D (nx10793), .CLK (clk), .R (rst)) ;
    mux21_ni ix10794 (.Y (nx10793), .A0 (camera_module_cache_ram_148__3), .A1 (
             nx35312), .S0 (nx34818)) ;
    aoi22 ix30325 (.Y (nx30324), .A0 (camera_module_cache_ram_180__3), .A1 (
          nx36232), .B0 (camera_module_cache_ram_164__3), .B1 (nx36272)) ;
    dffr camera_module_cache_reg_ram_180__3 (.Q (camera_module_cache_ram_180__3)
         , .QB (\$dummy [1384]), .D (nx10773), .CLK (clk), .R (rst)) ;
    mux21_ni ix10774 (.Y (nx10773), .A0 (camera_module_cache_ram_180__3), .A1 (
             nx35312), .S0 (nx34810)) ;
    dffr camera_module_cache_reg_ram_164__3 (.Q (camera_module_cache_ram_164__3)
         , .QB (\$dummy [1385]), .D (nx10783), .CLK (clk), .R (rst)) ;
    mux21_ni ix10784 (.Y (nx10783), .A0 (camera_module_cache_ram_164__3), .A1 (
             nx35312), .S0 (nx34814)) ;
    aoi22 ix30333 (.Y (nx30332), .A0 (camera_module_cache_ram_196__3), .A1 (
          nx36312), .B0 (camera_module_cache_ram_212__3), .B1 (nx36352)) ;
    dffr camera_module_cache_reg_ram_196__3 (.Q (camera_module_cache_ram_196__3)
         , .QB (\$dummy [1386]), .D (nx10763), .CLK (clk), .R (rst)) ;
    mux21_ni ix10764 (.Y (nx10763), .A0 (camera_module_cache_ram_196__3), .A1 (
             nx35312), .S0 (nx34806)) ;
    dffr camera_module_cache_reg_ram_212__3 (.Q (camera_module_cache_ram_212__3)
         , .QB (\$dummy [1387]), .D (nx10753), .CLK (clk), .R (rst)) ;
    mux21_ni ix10754 (.Y (nx10753), .A0 (camera_module_cache_ram_212__3), .A1 (
             nx35314), .S0 (nx34802)) ;
    aoi22 ix30341 (.Y (nx30340), .A0 (camera_module_cache_ram_228__3), .A1 (
          nx36392), .B0 (camera_module_cache_ram_244__3), .B1 (nx36432)) ;
    dffr camera_module_cache_reg_ram_228__3 (.Q (camera_module_cache_ram_228__3)
         , .QB (\$dummy [1388]), .D (nx10743), .CLK (clk), .R (rst)) ;
    mux21_ni ix10744 (.Y (nx10743), .A0 (camera_module_cache_ram_228__3), .A1 (
             nx35314), .S0 (nx34798)) ;
    dffr camera_module_cache_reg_ram_244__3 (.Q (camera_module_cache_ram_244__3)
         , .QB (\$dummy [1389]), .D (nx10733), .CLK (clk), .R (rst)) ;
    mux21_ni ix10734 (.Y (nx10733), .A0 (camera_module_cache_ram_244__3), .A1 (
             nx35314), .S0 (nx34794)) ;
    oai21 ix30349 (.Y (nx30348), .A0 (nx13440), .A1 (nx13362), .B0 (nx36468)) ;
    nand04 ix13441 (.Y (nx13440), .A0 (nx30351), .A1 (nx30359), .A2 (nx30367), .A3 (
           nx30375)) ;
    aoi22 ix30352 (.Y (nx30351), .A0 (camera_module_cache_ram_5__3), .A1 (
          nx35832), .B0 (camera_module_cache_ram_21__3), .B1 (nx35872)) ;
    dffr camera_module_cache_reg_ram_5__3 (.Q (camera_module_cache_ram_5__3), .QB (
         \$dummy [1390]), .D (nx10723), .CLK (clk), .R (rst)) ;
    mux21_ni ix10724 (.Y (nx10723), .A0 (camera_module_cache_ram_5__3), .A1 (
             nx35314), .S0 (nx34784)) ;
    dffr camera_module_cache_reg_ram_21__3 (.Q (camera_module_cache_ram_21__3), 
         .QB (\$dummy [1391]), .D (nx10713), .CLK (clk), .R (rst)) ;
    mux21_ni ix10714 (.Y (nx10713), .A0 (camera_module_cache_ram_21__3), .A1 (
             nx35314), .S0 (nx34780)) ;
    aoi22 ix30360 (.Y (nx30359), .A0 (camera_module_cache_ram_37__3), .A1 (
          nx35912), .B0 (camera_module_cache_ram_53__3), .B1 (nx35952)) ;
    dffr camera_module_cache_reg_ram_37__3 (.Q (camera_module_cache_ram_37__3), 
         .QB (\$dummy [1392]), .D (nx10703), .CLK (clk), .R (rst)) ;
    mux21_ni ix10704 (.Y (nx10703), .A0 (camera_module_cache_ram_37__3), .A1 (
             nx35314), .S0 (nx34776)) ;
    dffr camera_module_cache_reg_ram_53__3 (.Q (camera_module_cache_ram_53__3), 
         .QB (\$dummy [1393]), .D (nx10693), .CLK (clk), .R (rst)) ;
    mux21_ni ix10694 (.Y (nx10693), .A0 (camera_module_cache_ram_53__3), .A1 (
             nx35314), .S0 (nx34772)) ;
    aoi22 ix30368 (.Y (nx30367), .A0 (camera_module_cache_ram_69__3), .A1 (
          nx35992), .B0 (camera_module_cache_ram_85__3), .B1 (nx36032)) ;
    dffr camera_module_cache_reg_ram_69__3 (.Q (camera_module_cache_ram_69__3), 
         .QB (\$dummy [1394]), .D (nx10683), .CLK (clk), .R (rst)) ;
    mux21_ni ix10684 (.Y (nx10683), .A0 (camera_module_cache_ram_69__3), .A1 (
             nx35316), .S0 (nx34768)) ;
    dffr camera_module_cache_reg_ram_85__3 (.Q (camera_module_cache_ram_85__3), 
         .QB (\$dummy [1395]), .D (nx10673), .CLK (clk), .R (rst)) ;
    mux21_ni ix10674 (.Y (nx10673), .A0 (camera_module_cache_ram_85__3), .A1 (
             nx35316), .S0 (nx34764)) ;
    aoi22 ix30376 (.Y (nx30375), .A0 (camera_module_cache_ram_117__3), .A1 (
          nx36072), .B0 (camera_module_cache_ram_101__3), .B1 (nx36112)) ;
    dffr camera_module_cache_reg_ram_117__3 (.Q (camera_module_cache_ram_117__3)
         , .QB (\$dummy [1396]), .D (nx10653), .CLK (clk), .R (rst)) ;
    mux21_ni ix10654 (.Y (nx10653), .A0 (camera_module_cache_ram_117__3), .A1 (
             nx35316), .S0 (nx34756)) ;
    dffr camera_module_cache_reg_ram_101__3 (.Q (camera_module_cache_ram_101__3)
         , .QB (\$dummy [1397]), .D (nx10663), .CLK (clk), .R (rst)) ;
    mux21_ni ix10664 (.Y (nx10663), .A0 (camera_module_cache_ram_101__3), .A1 (
             nx35316), .S0 (nx34760)) ;
    nand04 ix13363 (.Y (nx13362), .A0 (nx30384), .A1 (nx30392), .A2 (nx30400), .A3 (
           nx30408)) ;
    aoi22 ix30385 (.Y (nx30384), .A0 (camera_module_cache_ram_133__3), .A1 (
          nx36152), .B0 (camera_module_cache_ram_149__3), .B1 (nx36192)) ;
    dffr camera_module_cache_reg_ram_133__3 (.Q (camera_module_cache_ram_133__3)
         , .QB (\$dummy [1398]), .D (nx10643), .CLK (clk), .R (rst)) ;
    mux21_ni ix10644 (.Y (nx10643), .A0 (camera_module_cache_ram_133__3), .A1 (
             nx35316), .S0 (nx34752)) ;
    dffr camera_module_cache_reg_ram_149__3 (.Q (camera_module_cache_ram_149__3)
         , .QB (\$dummy [1399]), .D (nx10633), .CLK (clk), .R (rst)) ;
    mux21_ni ix10634 (.Y (nx10633), .A0 (camera_module_cache_ram_149__3), .A1 (
             nx35316), .S0 (nx34748)) ;
    aoi22 ix30393 (.Y (nx30392), .A0 (camera_module_cache_ram_181__3), .A1 (
          nx36232), .B0 (camera_module_cache_ram_165__3), .B1 (nx36272)) ;
    dffr camera_module_cache_reg_ram_181__3 (.Q (camera_module_cache_ram_181__3)
         , .QB (\$dummy [1400]), .D (nx10613), .CLK (clk), .R (rst)) ;
    mux21_ni ix10614 (.Y (nx10613), .A0 (camera_module_cache_ram_181__3), .A1 (
             nx35316), .S0 (nx34740)) ;
    dffr camera_module_cache_reg_ram_165__3 (.Q (camera_module_cache_ram_165__3)
         , .QB (\$dummy [1401]), .D (nx10623), .CLK (clk), .R (rst)) ;
    mux21_ni ix10624 (.Y (nx10623), .A0 (camera_module_cache_ram_165__3), .A1 (
             nx35318), .S0 (nx34744)) ;
    aoi22 ix30401 (.Y (nx30400), .A0 (camera_module_cache_ram_197__3), .A1 (
          nx36312), .B0 (camera_module_cache_ram_213__3), .B1 (nx36352)) ;
    dffr camera_module_cache_reg_ram_197__3 (.Q (camera_module_cache_ram_197__3)
         , .QB (\$dummy [1402]), .D (nx10603), .CLK (clk), .R (rst)) ;
    mux21_ni ix10604 (.Y (nx10603), .A0 (camera_module_cache_ram_197__3), .A1 (
             nx35318), .S0 (nx34736)) ;
    dffr camera_module_cache_reg_ram_213__3 (.Q (camera_module_cache_ram_213__3)
         , .QB (\$dummy [1403]), .D (nx10593), .CLK (clk), .R (rst)) ;
    mux21_ni ix10594 (.Y (nx10593), .A0 (camera_module_cache_ram_213__3), .A1 (
             nx35318), .S0 (nx34732)) ;
    aoi22 ix30409 (.Y (nx30408), .A0 (camera_module_cache_ram_229__3), .A1 (
          nx36392), .B0 (camera_module_cache_ram_245__3), .B1 (nx36432)) ;
    dffr camera_module_cache_reg_ram_229__3 (.Q (camera_module_cache_ram_229__3)
         , .QB (\$dummy [1404]), .D (nx10583), .CLK (clk), .R (rst)) ;
    mux21_ni ix10584 (.Y (nx10583), .A0 (camera_module_cache_ram_229__3), .A1 (
             nx35318), .S0 (nx34728)) ;
    dffr camera_module_cache_reg_ram_245__3 (.Q (camera_module_cache_ram_245__3)
         , .QB (\$dummy [1405]), .D (nx10573), .CLK (clk), .R (rst)) ;
    mux21_ni ix10574 (.Y (nx10573), .A0 (camera_module_cache_ram_245__3), .A1 (
             nx35318), .S0 (nx34724)) ;
    oai21 ix30417 (.Y (nx30416), .A0 (nx13276), .A1 (nx13198), .B0 (nx36472)) ;
    nand04 ix13277 (.Y (nx13276), .A0 (nx30419), .A1 (nx30427), .A2 (nx30435), .A3 (
           nx30443)) ;
    aoi22 ix30420 (.Y (nx30419), .A0 (camera_module_cache_ram_6__3), .A1 (
          nx35832), .B0 (camera_module_cache_ram_22__3), .B1 (nx35872)) ;
    dffr camera_module_cache_reg_ram_6__3 (.Q (camera_module_cache_ram_6__3), .QB (
         \$dummy [1406]), .D (nx10563), .CLK (clk), .R (rst)) ;
    mux21_ni ix10564 (.Y (nx10563), .A0 (camera_module_cache_ram_6__3), .A1 (
             nx35318), .S0 (nx34714)) ;
    dffr camera_module_cache_reg_ram_22__3 (.Q (camera_module_cache_ram_22__3), 
         .QB (\$dummy [1407]), .D (nx10553), .CLK (clk), .R (rst)) ;
    mux21_ni ix10554 (.Y (nx10553), .A0 (camera_module_cache_ram_22__3), .A1 (
             nx35318), .S0 (nx34710)) ;
    aoi22 ix30428 (.Y (nx30427), .A0 (camera_module_cache_ram_38__3), .A1 (
          nx35912), .B0 (camera_module_cache_ram_54__3), .B1 (nx35952)) ;
    dffr camera_module_cache_reg_ram_38__3 (.Q (camera_module_cache_ram_38__3), 
         .QB (\$dummy [1408]), .D (nx10543), .CLK (clk), .R (rst)) ;
    mux21_ni ix10544 (.Y (nx10543), .A0 (camera_module_cache_ram_38__3), .A1 (
             nx35320), .S0 (nx34706)) ;
    dffr camera_module_cache_reg_ram_54__3 (.Q (camera_module_cache_ram_54__3), 
         .QB (\$dummy [1409]), .D (nx10533), .CLK (clk), .R (rst)) ;
    mux21_ni ix10534 (.Y (nx10533), .A0 (camera_module_cache_ram_54__3), .A1 (
             nx35320), .S0 (nx34702)) ;
    aoi22 ix30436 (.Y (nx30435), .A0 (camera_module_cache_ram_70__3), .A1 (
          nx35992), .B0 (camera_module_cache_ram_86__3), .B1 (nx36032)) ;
    dffr camera_module_cache_reg_ram_70__3 (.Q (camera_module_cache_ram_70__3), 
         .QB (\$dummy [1410]), .D (nx10523), .CLK (clk), .R (rst)) ;
    mux21_ni ix10524 (.Y (nx10523), .A0 (camera_module_cache_ram_70__3), .A1 (
             nx35320), .S0 (nx34698)) ;
    dffr camera_module_cache_reg_ram_86__3 (.Q (camera_module_cache_ram_86__3), 
         .QB (\$dummy [1411]), .D (nx10513), .CLK (clk), .R (rst)) ;
    mux21_ni ix10514 (.Y (nx10513), .A0 (camera_module_cache_ram_86__3), .A1 (
             nx35320), .S0 (nx34694)) ;
    aoi22 ix30444 (.Y (nx30443), .A0 (camera_module_cache_ram_118__3), .A1 (
          nx36072), .B0 (camera_module_cache_ram_102__3), .B1 (nx36112)) ;
    dffr camera_module_cache_reg_ram_118__3 (.Q (camera_module_cache_ram_118__3)
         , .QB (\$dummy [1412]), .D (nx10493), .CLK (clk), .R (rst)) ;
    mux21_ni ix10494 (.Y (nx10493), .A0 (camera_module_cache_ram_118__3), .A1 (
             nx35320), .S0 (nx34686)) ;
    dffr camera_module_cache_reg_ram_102__3 (.Q (camera_module_cache_ram_102__3)
         , .QB (\$dummy [1413]), .D (nx10503), .CLK (clk), .R (rst)) ;
    mux21_ni ix10504 (.Y (nx10503), .A0 (camera_module_cache_ram_102__3), .A1 (
             nx35320), .S0 (nx34690)) ;
    nand04 ix13199 (.Y (nx13198), .A0 (nx30452), .A1 (nx30460), .A2 (nx30468), .A3 (
           nx30476)) ;
    aoi22 ix30453 (.Y (nx30452), .A0 (camera_module_cache_ram_134__3), .A1 (
          nx36152), .B0 (camera_module_cache_ram_150__3), .B1 (nx36192)) ;
    dffr camera_module_cache_reg_ram_134__3 (.Q (camera_module_cache_ram_134__3)
         , .QB (\$dummy [1414]), .D (nx10483), .CLK (clk), .R (rst)) ;
    mux21_ni ix10484 (.Y (nx10483), .A0 (camera_module_cache_ram_134__3), .A1 (
             nx35320), .S0 (nx34682)) ;
    dffr camera_module_cache_reg_ram_150__3 (.Q (camera_module_cache_ram_150__3)
         , .QB (\$dummy [1415]), .D (nx10473), .CLK (clk), .R (rst)) ;
    mux21_ni ix10474 (.Y (nx10473), .A0 (camera_module_cache_ram_150__3), .A1 (
             nx35322), .S0 (nx34678)) ;
    aoi22 ix30461 (.Y (nx30460), .A0 (camera_module_cache_ram_182__3), .A1 (
          nx36232), .B0 (camera_module_cache_ram_166__3), .B1 (nx36272)) ;
    dffr camera_module_cache_reg_ram_182__3 (.Q (camera_module_cache_ram_182__3)
         , .QB (\$dummy [1416]), .D (nx10453), .CLK (clk), .R (rst)) ;
    mux21_ni ix10454 (.Y (nx10453), .A0 (camera_module_cache_ram_182__3), .A1 (
             nx35322), .S0 (nx34670)) ;
    dffr camera_module_cache_reg_ram_166__3 (.Q (camera_module_cache_ram_166__3)
         , .QB (\$dummy [1417]), .D (nx10463), .CLK (clk), .R (rst)) ;
    mux21_ni ix10464 (.Y (nx10463), .A0 (camera_module_cache_ram_166__3), .A1 (
             nx35322), .S0 (nx34674)) ;
    aoi22 ix30469 (.Y (nx30468), .A0 (camera_module_cache_ram_198__3), .A1 (
          nx36312), .B0 (camera_module_cache_ram_214__3), .B1 (nx36352)) ;
    dffr camera_module_cache_reg_ram_198__3 (.Q (camera_module_cache_ram_198__3)
         , .QB (\$dummy [1418]), .D (nx10443), .CLK (clk), .R (rst)) ;
    mux21_ni ix10444 (.Y (nx10443), .A0 (camera_module_cache_ram_198__3), .A1 (
             nx35322), .S0 (nx34666)) ;
    dffr camera_module_cache_reg_ram_214__3 (.Q (camera_module_cache_ram_214__3)
         , .QB (\$dummy [1419]), .D (nx10433), .CLK (clk), .R (rst)) ;
    mux21_ni ix10434 (.Y (nx10433), .A0 (camera_module_cache_ram_214__3), .A1 (
             nx35322), .S0 (nx34662)) ;
    aoi22 ix30477 (.Y (nx30476), .A0 (camera_module_cache_ram_230__3), .A1 (
          nx36392), .B0 (camera_module_cache_ram_246__3), .B1 (nx36432)) ;
    dffr camera_module_cache_reg_ram_230__3 (.Q (camera_module_cache_ram_230__3)
         , .QB (\$dummy [1420]), .D (nx10423), .CLK (clk), .R (rst)) ;
    mux21_ni ix10424 (.Y (nx10423), .A0 (camera_module_cache_ram_230__3), .A1 (
             nx35322), .S0 (nx34658)) ;
    dffr camera_module_cache_reg_ram_246__3 (.Q (camera_module_cache_ram_246__3)
         , .QB (\$dummy [1421]), .D (nx10413), .CLK (clk), .R (rst)) ;
    mux21_ni ix10414 (.Y (nx10413), .A0 (camera_module_cache_ram_246__3), .A1 (
             nx35322), .S0 (nx34654)) ;
    oai21 ix30485 (.Y (nx30484), .A0 (nx13114), .A1 (nx13036), .B0 (nx36476)) ;
    nand04 ix13115 (.Y (nx13114), .A0 (nx30487), .A1 (nx30495), .A2 (nx30503), .A3 (
           nx30511)) ;
    aoi22 ix30488 (.Y (nx30487), .A0 (camera_module_cache_ram_7__3), .A1 (
          nx35834), .B0 (camera_module_cache_ram_23__3), .B1 (nx35874)) ;
    dffr camera_module_cache_reg_ram_7__3 (.Q (camera_module_cache_ram_7__3), .QB (
         \$dummy [1422]), .D (nx10403), .CLK (clk), .R (rst)) ;
    mux21_ni ix10404 (.Y (nx10403), .A0 (camera_module_cache_ram_7__3), .A1 (
             nx35324), .S0 (nx34644)) ;
    dffr camera_module_cache_reg_ram_23__3 (.Q (camera_module_cache_ram_23__3), 
         .QB (\$dummy [1423]), .D (nx10393), .CLK (clk), .R (rst)) ;
    mux21_ni ix10394 (.Y (nx10393), .A0 (camera_module_cache_ram_23__3), .A1 (
             nx35324), .S0 (nx34640)) ;
    aoi22 ix30496 (.Y (nx30495), .A0 (camera_module_cache_ram_39__3), .A1 (
          nx35914), .B0 (camera_module_cache_ram_55__3), .B1 (nx35954)) ;
    dffr camera_module_cache_reg_ram_39__3 (.Q (camera_module_cache_ram_39__3), 
         .QB (\$dummy [1424]), .D (nx10383), .CLK (clk), .R (rst)) ;
    mux21_ni ix10384 (.Y (nx10383), .A0 (camera_module_cache_ram_39__3), .A1 (
             nx35324), .S0 (nx34636)) ;
    dffr camera_module_cache_reg_ram_55__3 (.Q (camera_module_cache_ram_55__3), 
         .QB (\$dummy [1425]), .D (nx10373), .CLK (clk), .R (rst)) ;
    mux21_ni ix10374 (.Y (nx10373), .A0 (camera_module_cache_ram_55__3), .A1 (
             nx35324), .S0 (nx34632)) ;
    aoi22 ix30504 (.Y (nx30503), .A0 (camera_module_cache_ram_71__3), .A1 (
          nx35994), .B0 (camera_module_cache_ram_87__3), .B1 (nx36034)) ;
    dffr camera_module_cache_reg_ram_71__3 (.Q (camera_module_cache_ram_71__3), 
         .QB (\$dummy [1426]), .D (nx10363), .CLK (clk), .R (rst)) ;
    mux21_ni ix10364 (.Y (nx10363), .A0 (camera_module_cache_ram_71__3), .A1 (
             nx35324), .S0 (nx34628)) ;
    dffr camera_module_cache_reg_ram_87__3 (.Q (camera_module_cache_ram_87__3), 
         .QB (\$dummy [1427]), .D (nx10353), .CLK (clk), .R (rst)) ;
    mux21_ni ix10354 (.Y (nx10353), .A0 (camera_module_cache_ram_87__3), .A1 (
             nx35324), .S0 (nx34624)) ;
    aoi22 ix30512 (.Y (nx30511), .A0 (camera_module_cache_ram_119__3), .A1 (
          nx36074), .B0 (camera_module_cache_ram_103__3), .B1 (nx36114)) ;
    dffr camera_module_cache_reg_ram_119__3 (.Q (camera_module_cache_ram_119__3)
         , .QB (\$dummy [1428]), .D (nx10333), .CLK (clk), .R (rst)) ;
    mux21_ni ix10334 (.Y (nx10333), .A0 (camera_module_cache_ram_119__3), .A1 (
             nx35324), .S0 (nx34616)) ;
    dffr camera_module_cache_reg_ram_103__3 (.Q (camera_module_cache_ram_103__3)
         , .QB (\$dummy [1429]), .D (nx10343), .CLK (clk), .R (rst)) ;
    mux21_ni ix10344 (.Y (nx10343), .A0 (camera_module_cache_ram_103__3), .A1 (
             nx35326), .S0 (nx34620)) ;
    nand04 ix13037 (.Y (nx13036), .A0 (nx30520), .A1 (nx30528), .A2 (nx30536), .A3 (
           nx30544)) ;
    aoi22 ix30521 (.Y (nx30520), .A0 (camera_module_cache_ram_135__3), .A1 (
          nx36154), .B0 (camera_module_cache_ram_151__3), .B1 (nx36194)) ;
    dffr camera_module_cache_reg_ram_135__3 (.Q (camera_module_cache_ram_135__3)
         , .QB (\$dummy [1430]), .D (nx10323), .CLK (clk), .R (rst)) ;
    mux21_ni ix10324 (.Y (nx10323), .A0 (camera_module_cache_ram_135__3), .A1 (
             nx35326), .S0 (nx34612)) ;
    dffr camera_module_cache_reg_ram_151__3 (.Q (camera_module_cache_ram_151__3)
         , .QB (\$dummy [1431]), .D (nx10313), .CLK (clk), .R (rst)) ;
    mux21_ni ix10314 (.Y (nx10313), .A0 (camera_module_cache_ram_151__3), .A1 (
             nx35326), .S0 (nx34608)) ;
    aoi22 ix30529 (.Y (nx30528), .A0 (camera_module_cache_ram_183__3), .A1 (
          nx36234), .B0 (camera_module_cache_ram_167__3), .B1 (nx36274)) ;
    dffr camera_module_cache_reg_ram_183__3 (.Q (camera_module_cache_ram_183__3)
         , .QB (\$dummy [1432]), .D (nx10293), .CLK (clk), .R (rst)) ;
    mux21_ni ix10294 (.Y (nx10293), .A0 (camera_module_cache_ram_183__3), .A1 (
             nx35326), .S0 (nx34600)) ;
    dffr camera_module_cache_reg_ram_167__3 (.Q (camera_module_cache_ram_167__3)
         , .QB (\$dummy [1433]), .D (nx10303), .CLK (clk), .R (rst)) ;
    mux21_ni ix10304 (.Y (nx10303), .A0 (camera_module_cache_ram_167__3), .A1 (
             nx35326), .S0 (nx34604)) ;
    aoi22 ix30537 (.Y (nx30536), .A0 (camera_module_cache_ram_199__3), .A1 (
          nx36314), .B0 (camera_module_cache_ram_215__3), .B1 (nx36354)) ;
    dffr camera_module_cache_reg_ram_199__3 (.Q (camera_module_cache_ram_199__3)
         , .QB (\$dummy [1434]), .D (nx10283), .CLK (clk), .R (rst)) ;
    mux21_ni ix10284 (.Y (nx10283), .A0 (camera_module_cache_ram_199__3), .A1 (
             nx35326), .S0 (nx34596)) ;
    dffr camera_module_cache_reg_ram_215__3 (.Q (camera_module_cache_ram_215__3)
         , .QB (\$dummy [1435]), .D (nx10273), .CLK (clk), .R (rst)) ;
    mux21_ni ix10274 (.Y (nx10273), .A0 (camera_module_cache_ram_215__3), .A1 (
             nx35326), .S0 (nx34592)) ;
    aoi22 ix30545 (.Y (nx30544), .A0 (camera_module_cache_ram_231__3), .A1 (
          nx36394), .B0 (camera_module_cache_ram_247__3), .B1 (nx36434)) ;
    dffr camera_module_cache_reg_ram_231__3 (.Q (camera_module_cache_ram_231__3)
         , .QB (\$dummy [1436]), .D (nx10263), .CLK (clk), .R (rst)) ;
    mux21_ni ix10264 (.Y (nx10263), .A0 (camera_module_cache_ram_231__3), .A1 (
             nx35328), .S0 (nx34588)) ;
    dffr camera_module_cache_reg_ram_247__3 (.Q (camera_module_cache_ram_247__3)
         , .QB (\$dummy [1437]), .D (nx10253), .CLK (clk), .R (rst)) ;
    mux21_ni ix10254 (.Y (nx10253), .A0 (camera_module_cache_ram_247__3), .A1 (
             nx35328), .S0 (nx34584)) ;
    nand04 ix12957 (.Y (nx12956), .A0 (nx30553), .A1 (nx30621), .A2 (nx30689), .A3 (
           nx30757)) ;
    oai21 ix30554 (.Y (nx30553), .A0 (nx12946), .A1 (nx12868), .B0 (nx36480)) ;
    nand04 ix12947 (.Y (nx12946), .A0 (nx30556), .A1 (nx30564), .A2 (nx30572), .A3 (
           nx30580)) ;
    aoi22 ix30557 (.Y (nx30556), .A0 (camera_module_cache_ram_8__3), .A1 (
          nx35834), .B0 (camera_module_cache_ram_24__3), .B1 (nx35874)) ;
    dffr camera_module_cache_reg_ram_8__3 (.Q (camera_module_cache_ram_8__3), .QB (
         \$dummy [1438]), .D (nx10243), .CLK (clk), .R (rst)) ;
    mux21_ni ix10244 (.Y (nx10243), .A0 (camera_module_cache_ram_8__3), .A1 (
             nx35328), .S0 (nx34574)) ;
    dffr camera_module_cache_reg_ram_24__3 (.Q (camera_module_cache_ram_24__3), 
         .QB (\$dummy [1439]), .D (nx10233), .CLK (clk), .R (rst)) ;
    mux21_ni ix10234 (.Y (nx10233), .A0 (camera_module_cache_ram_24__3), .A1 (
             nx35328), .S0 (nx34570)) ;
    aoi22 ix30565 (.Y (nx30564), .A0 (camera_module_cache_ram_40__3), .A1 (
          nx35914), .B0 (camera_module_cache_ram_56__3), .B1 (nx35954)) ;
    dffr camera_module_cache_reg_ram_40__3 (.Q (camera_module_cache_ram_40__3), 
         .QB (\$dummy [1440]), .D (nx10223), .CLK (clk), .R (rst)) ;
    mux21_ni ix10224 (.Y (nx10223), .A0 (camera_module_cache_ram_40__3), .A1 (
             nx35328), .S0 (nx34566)) ;
    dffr camera_module_cache_reg_ram_56__3 (.Q (camera_module_cache_ram_56__3), 
         .QB (\$dummy [1441]), .D (nx10213), .CLK (clk), .R (rst)) ;
    mux21_ni ix10214 (.Y (nx10213), .A0 (camera_module_cache_ram_56__3), .A1 (
             nx35328), .S0 (nx34562)) ;
    aoi22 ix30573 (.Y (nx30572), .A0 (camera_module_cache_ram_72__3), .A1 (
          nx35994), .B0 (camera_module_cache_ram_88__3), .B1 (nx36034)) ;
    dffr camera_module_cache_reg_ram_72__3 (.Q (camera_module_cache_ram_72__3), 
         .QB (\$dummy [1442]), .D (nx10203), .CLK (clk), .R (rst)) ;
    mux21_ni ix10204 (.Y (nx10203), .A0 (camera_module_cache_ram_72__3), .A1 (
             nx35328), .S0 (nx34558)) ;
    dffr camera_module_cache_reg_ram_88__3 (.Q (camera_module_cache_ram_88__3), 
         .QB (\$dummy [1443]), .D (nx10193), .CLK (clk), .R (rst)) ;
    mux21_ni ix10194 (.Y (nx10193), .A0 (camera_module_cache_ram_88__3), .A1 (
             nx35330), .S0 (nx34554)) ;
    aoi22 ix30581 (.Y (nx30580), .A0 (camera_module_cache_ram_120__3), .A1 (
          nx36074), .B0 (camera_module_cache_ram_104__3), .B1 (nx36114)) ;
    dffr camera_module_cache_reg_ram_120__3 (.Q (camera_module_cache_ram_120__3)
         , .QB (\$dummy [1444]), .D (nx10173), .CLK (clk), .R (rst)) ;
    mux21_ni ix10174 (.Y (nx10173), .A0 (camera_module_cache_ram_120__3), .A1 (
             nx35330), .S0 (nx34546)) ;
    dffr camera_module_cache_reg_ram_104__3 (.Q (camera_module_cache_ram_104__3)
         , .QB (\$dummy [1445]), .D (nx10183), .CLK (clk), .R (rst)) ;
    mux21_ni ix10184 (.Y (nx10183), .A0 (camera_module_cache_ram_104__3), .A1 (
             nx35330), .S0 (nx34550)) ;
    nand04 ix12869 (.Y (nx12868), .A0 (nx30589), .A1 (nx30597), .A2 (nx30605), .A3 (
           nx30613)) ;
    aoi22 ix30590 (.Y (nx30589), .A0 (camera_module_cache_ram_136__3), .A1 (
          nx36154), .B0 (camera_module_cache_ram_152__3), .B1 (nx36194)) ;
    dffr camera_module_cache_reg_ram_136__3 (.Q (camera_module_cache_ram_136__3)
         , .QB (\$dummy [1446]), .D (nx10163), .CLK (clk), .R (rst)) ;
    mux21_ni ix10164 (.Y (nx10163), .A0 (camera_module_cache_ram_136__3), .A1 (
             nx35330), .S0 (nx34542)) ;
    dffr camera_module_cache_reg_ram_152__3 (.Q (camera_module_cache_ram_152__3)
         , .QB (\$dummy [1447]), .D (nx10153), .CLK (clk), .R (rst)) ;
    mux21_ni ix10154 (.Y (nx10153), .A0 (camera_module_cache_ram_152__3), .A1 (
             nx35330), .S0 (nx34538)) ;
    aoi22 ix30598 (.Y (nx30597), .A0 (camera_module_cache_ram_184__3), .A1 (
          nx36234), .B0 (camera_module_cache_ram_168__3), .B1 (nx36274)) ;
    dffr camera_module_cache_reg_ram_184__3 (.Q (camera_module_cache_ram_184__3)
         , .QB (\$dummy [1448]), .D (nx10133), .CLK (clk), .R (rst)) ;
    mux21_ni ix10134 (.Y (nx10133), .A0 (camera_module_cache_ram_184__3), .A1 (
             nx35330), .S0 (nx34530)) ;
    dffr camera_module_cache_reg_ram_168__3 (.Q (camera_module_cache_ram_168__3)
         , .QB (\$dummy [1449]), .D (nx10143), .CLK (clk), .R (rst)) ;
    mux21_ni ix10144 (.Y (nx10143), .A0 (camera_module_cache_ram_168__3), .A1 (
             nx35330), .S0 (nx34534)) ;
    aoi22 ix30606 (.Y (nx30605), .A0 (camera_module_cache_ram_200__3), .A1 (
          nx36314), .B0 (camera_module_cache_ram_216__3), .B1 (nx36354)) ;
    dffr camera_module_cache_reg_ram_200__3 (.Q (camera_module_cache_ram_200__3)
         , .QB (\$dummy [1450]), .D (nx10123), .CLK (clk), .R (rst)) ;
    mux21_ni ix10124 (.Y (nx10123), .A0 (camera_module_cache_ram_200__3), .A1 (
             nx35332), .S0 (nx34526)) ;
    dffr camera_module_cache_reg_ram_216__3 (.Q (camera_module_cache_ram_216__3)
         , .QB (\$dummy [1451]), .D (nx10113), .CLK (clk), .R (rst)) ;
    mux21_ni ix10114 (.Y (nx10113), .A0 (camera_module_cache_ram_216__3), .A1 (
             nx35332), .S0 (nx34522)) ;
    aoi22 ix30614 (.Y (nx30613), .A0 (camera_module_cache_ram_232__3), .A1 (
          nx36394), .B0 (camera_module_cache_ram_248__3), .B1 (nx36434)) ;
    dffr camera_module_cache_reg_ram_232__3 (.Q (camera_module_cache_ram_232__3)
         , .QB (\$dummy [1452]), .D (nx10103), .CLK (clk), .R (rst)) ;
    mux21_ni ix10104 (.Y (nx10103), .A0 (camera_module_cache_ram_232__3), .A1 (
             nx35332), .S0 (nx34518)) ;
    dffr camera_module_cache_reg_ram_248__3 (.Q (camera_module_cache_ram_248__3)
         , .QB (\$dummy [1453]), .D (nx10093), .CLK (clk), .R (rst)) ;
    mux21_ni ix10094 (.Y (nx10093), .A0 (camera_module_cache_ram_248__3), .A1 (
             nx35332), .S0 (nx34514)) ;
    oai21 ix30622 (.Y (nx30621), .A0 (nx12784), .A1 (nx12706), .B0 (nx36484)) ;
    nand04 ix12785 (.Y (nx12784), .A0 (nx30624), .A1 (nx30632), .A2 (nx30640), .A3 (
           nx30648)) ;
    aoi22 ix30625 (.Y (nx30624), .A0 (camera_module_cache_ram_9__3), .A1 (
          nx35834), .B0 (camera_module_cache_ram_25__3), .B1 (nx35874)) ;
    dffr camera_module_cache_reg_ram_9__3 (.Q (camera_module_cache_ram_9__3), .QB (
         \$dummy [1454]), .D (nx10083), .CLK (clk), .R (rst)) ;
    mux21_ni ix10084 (.Y (nx10083), .A0 (camera_module_cache_ram_9__3), .A1 (
             nx35332), .S0 (nx34504)) ;
    dffr camera_module_cache_reg_ram_25__3 (.Q (camera_module_cache_ram_25__3), 
         .QB (\$dummy [1455]), .D (nx10073), .CLK (clk), .R (rst)) ;
    mux21_ni ix10074 (.Y (nx10073), .A0 (camera_module_cache_ram_25__3), .A1 (
             nx35332), .S0 (nx34500)) ;
    aoi22 ix30633 (.Y (nx30632), .A0 (camera_module_cache_ram_41__3), .A1 (
          nx35914), .B0 (camera_module_cache_ram_57__3), .B1 (nx35954)) ;
    dffr camera_module_cache_reg_ram_41__3 (.Q (camera_module_cache_ram_41__3), 
         .QB (\$dummy [1456]), .D (nx10063), .CLK (clk), .R (rst)) ;
    mux21_ni ix10064 (.Y (nx10063), .A0 (camera_module_cache_ram_41__3), .A1 (
             nx35332), .S0 (nx34496)) ;
    dffr camera_module_cache_reg_ram_57__3 (.Q (camera_module_cache_ram_57__3), 
         .QB (\$dummy [1457]), .D (nx10053), .CLK (clk), .R (rst)) ;
    mux21_ni ix10054 (.Y (nx10053), .A0 (camera_module_cache_ram_57__3), .A1 (
             nx35334), .S0 (nx34492)) ;
    aoi22 ix30641 (.Y (nx30640), .A0 (camera_module_cache_ram_73__3), .A1 (
          nx35994), .B0 (camera_module_cache_ram_89__3), .B1 (nx36034)) ;
    dffr camera_module_cache_reg_ram_73__3 (.Q (camera_module_cache_ram_73__3), 
         .QB (\$dummy [1458]), .D (nx10043), .CLK (clk), .R (rst)) ;
    mux21_ni ix10044 (.Y (nx10043), .A0 (camera_module_cache_ram_73__3), .A1 (
             nx35334), .S0 (nx34488)) ;
    dffr camera_module_cache_reg_ram_89__3 (.Q (camera_module_cache_ram_89__3), 
         .QB (\$dummy [1459]), .D (nx10033), .CLK (clk), .R (rst)) ;
    mux21_ni ix10034 (.Y (nx10033), .A0 (camera_module_cache_ram_89__3), .A1 (
             nx35334), .S0 (nx34484)) ;
    aoi22 ix30649 (.Y (nx30648), .A0 (camera_module_cache_ram_121__3), .A1 (
          nx36074), .B0 (camera_module_cache_ram_105__3), .B1 (nx36114)) ;
    dffr camera_module_cache_reg_ram_121__3 (.Q (camera_module_cache_ram_121__3)
         , .QB (\$dummy [1460]), .D (nx10013), .CLK (clk), .R (rst)) ;
    mux21_ni ix10014 (.Y (nx10013), .A0 (camera_module_cache_ram_121__3), .A1 (
             nx35334), .S0 (nx34476)) ;
    dffr camera_module_cache_reg_ram_105__3 (.Q (camera_module_cache_ram_105__3)
         , .QB (\$dummy [1461]), .D (nx10023), .CLK (clk), .R (rst)) ;
    mux21_ni ix10024 (.Y (nx10023), .A0 (camera_module_cache_ram_105__3), .A1 (
             nx35334), .S0 (nx34480)) ;
    nand04 ix12707 (.Y (nx12706), .A0 (nx30657), .A1 (nx30665), .A2 (nx30673), .A3 (
           nx30681)) ;
    aoi22 ix30658 (.Y (nx30657), .A0 (camera_module_cache_ram_137__3), .A1 (
          nx36154), .B0 (camera_module_cache_ram_153__3), .B1 (nx36194)) ;
    dffr camera_module_cache_reg_ram_137__3 (.Q (camera_module_cache_ram_137__3)
         , .QB (\$dummy [1462]), .D (nx10003), .CLK (clk), .R (rst)) ;
    mux21_ni ix10004 (.Y (nx10003), .A0 (camera_module_cache_ram_137__3), .A1 (
             nx35334), .S0 (nx34472)) ;
    dffr camera_module_cache_reg_ram_153__3 (.Q (camera_module_cache_ram_153__3)
         , .QB (\$dummy [1463]), .D (nx9993), .CLK (clk), .R (rst)) ;
    mux21_ni ix9994 (.Y (nx9993), .A0 (camera_module_cache_ram_153__3), .A1 (
             nx35334), .S0 (nx34468)) ;
    aoi22 ix30666 (.Y (nx30665), .A0 (camera_module_cache_ram_185__3), .A1 (
          nx36234), .B0 (camera_module_cache_ram_169__3), .B1 (nx36274)) ;
    dffr camera_module_cache_reg_ram_185__3 (.Q (camera_module_cache_ram_185__3)
         , .QB (\$dummy [1464]), .D (nx9973), .CLK (clk), .R (rst)) ;
    mux21_ni ix9974 (.Y (nx9973), .A0 (camera_module_cache_ram_185__3), .A1 (
             nx35336), .S0 (nx34460)) ;
    dffr camera_module_cache_reg_ram_169__3 (.Q (camera_module_cache_ram_169__3)
         , .QB (\$dummy [1465]), .D (nx9983), .CLK (clk), .R (rst)) ;
    mux21_ni ix9984 (.Y (nx9983), .A0 (camera_module_cache_ram_169__3), .A1 (
             nx35336), .S0 (nx34464)) ;
    aoi22 ix30674 (.Y (nx30673), .A0 (camera_module_cache_ram_201__3), .A1 (
          nx36314), .B0 (camera_module_cache_ram_217__3), .B1 (nx36354)) ;
    dffr camera_module_cache_reg_ram_201__3 (.Q (camera_module_cache_ram_201__3)
         , .QB (\$dummy [1466]), .D (nx9963), .CLK (clk), .R (rst)) ;
    mux21_ni ix9964 (.Y (nx9963), .A0 (camera_module_cache_ram_201__3), .A1 (
             nx35336), .S0 (nx34456)) ;
    dffr camera_module_cache_reg_ram_217__3 (.Q (camera_module_cache_ram_217__3)
         , .QB (\$dummy [1467]), .D (nx9953), .CLK (clk), .R (rst)) ;
    mux21_ni ix9954 (.Y (nx9953), .A0 (camera_module_cache_ram_217__3), .A1 (
             nx35336), .S0 (nx34452)) ;
    aoi22 ix30682 (.Y (nx30681), .A0 (camera_module_cache_ram_233__3), .A1 (
          nx36394), .B0 (camera_module_cache_ram_249__3), .B1 (nx36434)) ;
    dffr camera_module_cache_reg_ram_233__3 (.Q (camera_module_cache_ram_233__3)
         , .QB (\$dummy [1468]), .D (nx9943), .CLK (clk), .R (rst)) ;
    mux21_ni ix9944 (.Y (nx9943), .A0 (camera_module_cache_ram_233__3), .A1 (
             nx35336), .S0 (nx34448)) ;
    dffr camera_module_cache_reg_ram_249__3 (.Q (camera_module_cache_ram_249__3)
         , .QB (\$dummy [1469]), .D (nx9933), .CLK (clk), .R (rst)) ;
    mux21_ni ix9934 (.Y (nx9933), .A0 (camera_module_cache_ram_249__3), .A1 (
             nx35336), .S0 (nx34444)) ;
    oai21 ix30690 (.Y (nx30689), .A0 (nx12620), .A1 (nx12542), .B0 (nx36488)) ;
    nand04 ix12621 (.Y (nx12620), .A0 (nx30692), .A1 (nx30700), .A2 (nx30708), .A3 (
           nx30716)) ;
    aoi22 ix30693 (.Y (nx30692), .A0 (camera_module_cache_ram_10__3), .A1 (
          nx35834), .B0 (camera_module_cache_ram_26__3), .B1 (nx35874)) ;
    dffr camera_module_cache_reg_ram_10__3 (.Q (camera_module_cache_ram_10__3), 
         .QB (\$dummy [1470]), .D (nx9923), .CLK (clk), .R (rst)) ;
    mux21_ni ix9924 (.Y (nx9923), .A0 (camera_module_cache_ram_10__3), .A1 (
             nx35336), .S0 (nx34434)) ;
    dffr camera_module_cache_reg_ram_26__3 (.Q (camera_module_cache_ram_26__3), 
         .QB (\$dummy [1471]), .D (nx9913), .CLK (clk), .R (rst)) ;
    mux21_ni ix9914 (.Y (nx9913), .A0 (camera_module_cache_ram_26__3), .A1 (
             nx35338), .S0 (nx34430)) ;
    aoi22 ix30701 (.Y (nx30700), .A0 (camera_module_cache_ram_42__3), .A1 (
          nx35914), .B0 (camera_module_cache_ram_58__3), .B1 (nx35954)) ;
    dffr camera_module_cache_reg_ram_42__3 (.Q (camera_module_cache_ram_42__3), 
         .QB (\$dummy [1472]), .D (nx9903), .CLK (clk), .R (rst)) ;
    mux21_ni ix9904 (.Y (nx9903), .A0 (camera_module_cache_ram_42__3), .A1 (
             nx35338), .S0 (nx34426)) ;
    dffr camera_module_cache_reg_ram_58__3 (.Q (camera_module_cache_ram_58__3), 
         .QB (\$dummy [1473]), .D (nx9893), .CLK (clk), .R (rst)) ;
    mux21_ni ix9894 (.Y (nx9893), .A0 (camera_module_cache_ram_58__3), .A1 (
             nx35338), .S0 (nx34422)) ;
    aoi22 ix30709 (.Y (nx30708), .A0 (camera_module_cache_ram_74__3), .A1 (
          nx35994), .B0 (camera_module_cache_ram_90__3), .B1 (nx36034)) ;
    dffr camera_module_cache_reg_ram_74__3 (.Q (camera_module_cache_ram_74__3), 
         .QB (\$dummy [1474]), .D (nx9883), .CLK (clk), .R (rst)) ;
    mux21_ni ix9884 (.Y (nx9883), .A0 (camera_module_cache_ram_74__3), .A1 (
             nx35338), .S0 (nx34418)) ;
    dffr camera_module_cache_reg_ram_90__3 (.Q (camera_module_cache_ram_90__3), 
         .QB (\$dummy [1475]), .D (nx9873), .CLK (clk), .R (rst)) ;
    mux21_ni ix9874 (.Y (nx9873), .A0 (camera_module_cache_ram_90__3), .A1 (
             nx35338), .S0 (nx34414)) ;
    aoi22 ix30717 (.Y (nx30716), .A0 (camera_module_cache_ram_122__3), .A1 (
          nx36074), .B0 (camera_module_cache_ram_106__3), .B1 (nx36114)) ;
    dffr camera_module_cache_reg_ram_122__3 (.Q (camera_module_cache_ram_122__3)
         , .QB (\$dummy [1476]), .D (nx9853), .CLK (clk), .R (rst)) ;
    mux21_ni ix9854 (.Y (nx9853), .A0 (camera_module_cache_ram_122__3), .A1 (
             nx35338), .S0 (nx34406)) ;
    dffr camera_module_cache_reg_ram_106__3 (.Q (camera_module_cache_ram_106__3)
         , .QB (\$dummy [1477]), .D (nx9863), .CLK (clk), .R (rst)) ;
    mux21_ni ix9864 (.Y (nx9863), .A0 (camera_module_cache_ram_106__3), .A1 (
             nx35338), .S0 (nx34410)) ;
    nand04 ix12543 (.Y (nx12542), .A0 (nx30725), .A1 (nx30733), .A2 (nx30741), .A3 (
           nx30749)) ;
    aoi22 ix30726 (.Y (nx30725), .A0 (camera_module_cache_ram_138__3), .A1 (
          nx36154), .B0 (camera_module_cache_ram_154__3), .B1 (nx36194)) ;
    dffr camera_module_cache_reg_ram_138__3 (.Q (camera_module_cache_ram_138__3)
         , .QB (\$dummy [1478]), .D (nx9843), .CLK (clk), .R (rst)) ;
    mux21_ni ix9844 (.Y (nx9843), .A0 (camera_module_cache_ram_138__3), .A1 (
             nx35340), .S0 (nx34402)) ;
    dffr camera_module_cache_reg_ram_154__3 (.Q (camera_module_cache_ram_154__3)
         , .QB (\$dummy [1479]), .D (nx9833), .CLK (clk), .R (rst)) ;
    mux21_ni ix9834 (.Y (nx9833), .A0 (camera_module_cache_ram_154__3), .A1 (
             nx35340), .S0 (nx34398)) ;
    aoi22 ix30734 (.Y (nx30733), .A0 (camera_module_cache_ram_186__3), .A1 (
          nx36234), .B0 (camera_module_cache_ram_170__3), .B1 (nx36274)) ;
    dffr camera_module_cache_reg_ram_186__3 (.Q (camera_module_cache_ram_186__3)
         , .QB (\$dummy [1480]), .D (nx9813), .CLK (clk), .R (rst)) ;
    mux21_ni ix9814 (.Y (nx9813), .A0 (camera_module_cache_ram_186__3), .A1 (
             nx35340), .S0 (nx34390)) ;
    dffr camera_module_cache_reg_ram_170__3 (.Q (camera_module_cache_ram_170__3)
         , .QB (\$dummy [1481]), .D (nx9823), .CLK (clk), .R (rst)) ;
    mux21_ni ix9824 (.Y (nx9823), .A0 (camera_module_cache_ram_170__3), .A1 (
             nx35340), .S0 (nx34394)) ;
    aoi22 ix30742 (.Y (nx30741), .A0 (camera_module_cache_ram_202__3), .A1 (
          nx36314), .B0 (camera_module_cache_ram_218__3), .B1 (nx36354)) ;
    dffr camera_module_cache_reg_ram_202__3 (.Q (camera_module_cache_ram_202__3)
         , .QB (\$dummy [1482]), .D (nx9803), .CLK (clk), .R (rst)) ;
    mux21_ni ix9804 (.Y (nx9803), .A0 (camera_module_cache_ram_202__3), .A1 (
             nx35340), .S0 (nx34386)) ;
    dffr camera_module_cache_reg_ram_218__3 (.Q (camera_module_cache_ram_218__3)
         , .QB (\$dummy [1483]), .D (nx9793), .CLK (clk), .R (rst)) ;
    mux21_ni ix9794 (.Y (nx9793), .A0 (camera_module_cache_ram_218__3), .A1 (
             nx35340), .S0 (nx34382)) ;
    aoi22 ix30750 (.Y (nx30749), .A0 (camera_module_cache_ram_234__3), .A1 (
          nx36394), .B0 (camera_module_cache_ram_250__3), .B1 (nx36434)) ;
    dffr camera_module_cache_reg_ram_234__3 (.Q (camera_module_cache_ram_234__3)
         , .QB (\$dummy [1484]), .D (nx9783), .CLK (clk), .R (rst)) ;
    mux21_ni ix9784 (.Y (nx9783), .A0 (camera_module_cache_ram_234__3), .A1 (
             nx35340), .S0 (nx34378)) ;
    dffr camera_module_cache_reg_ram_250__3 (.Q (camera_module_cache_ram_250__3)
         , .QB (\$dummy [1485]), .D (nx9773), .CLK (clk), .R (rst)) ;
    mux21_ni ix9774 (.Y (nx9773), .A0 (camera_module_cache_ram_250__3), .A1 (
             nx35342), .S0 (nx34374)) ;
    oai21 ix30758 (.Y (nx30757), .A0 (nx12458), .A1 (nx12380), .B0 (nx36492)) ;
    nand04 ix12459 (.Y (nx12458), .A0 (nx30760), .A1 (nx30768), .A2 (nx30776), .A3 (
           nx30784)) ;
    aoi22 ix30761 (.Y (nx30760), .A0 (camera_module_cache_ram_11__3), .A1 (
          nx35834), .B0 (camera_module_cache_ram_27__3), .B1 (nx35874)) ;
    dffr camera_module_cache_reg_ram_11__3 (.Q (camera_module_cache_ram_11__3), 
         .QB (\$dummy [1486]), .D (nx9763), .CLK (clk), .R (rst)) ;
    mux21_ni ix9764 (.Y (nx9763), .A0 (camera_module_cache_ram_11__3), .A1 (
             nx35342), .S0 (nx34364)) ;
    dffr camera_module_cache_reg_ram_27__3 (.Q (camera_module_cache_ram_27__3), 
         .QB (\$dummy [1487]), .D (nx9753), .CLK (clk), .R (rst)) ;
    mux21_ni ix9754 (.Y (nx9753), .A0 (camera_module_cache_ram_27__3), .A1 (
             nx35342), .S0 (nx34360)) ;
    aoi22 ix30769 (.Y (nx30768), .A0 (camera_module_cache_ram_43__3), .A1 (
          nx35914), .B0 (camera_module_cache_ram_59__3), .B1 (nx35954)) ;
    dffr camera_module_cache_reg_ram_43__3 (.Q (camera_module_cache_ram_43__3), 
         .QB (\$dummy [1488]), .D (nx9743), .CLK (clk), .R (rst)) ;
    mux21_ni ix9744 (.Y (nx9743), .A0 (camera_module_cache_ram_43__3), .A1 (
             nx35342), .S0 (nx34356)) ;
    dffr camera_module_cache_reg_ram_59__3 (.Q (camera_module_cache_ram_59__3), 
         .QB (\$dummy [1489]), .D (nx9733), .CLK (clk), .R (rst)) ;
    mux21_ni ix9734 (.Y (nx9733), .A0 (camera_module_cache_ram_59__3), .A1 (
             nx35342), .S0 (nx34352)) ;
    aoi22 ix30777 (.Y (nx30776), .A0 (camera_module_cache_ram_75__3), .A1 (
          nx35994), .B0 (camera_module_cache_ram_91__3), .B1 (nx36034)) ;
    dffr camera_module_cache_reg_ram_75__3 (.Q (camera_module_cache_ram_75__3), 
         .QB (\$dummy [1490]), .D (nx9723), .CLK (clk), .R (rst)) ;
    mux21_ni ix9724 (.Y (nx9723), .A0 (camera_module_cache_ram_75__3), .A1 (
             nx35342), .S0 (nx34348)) ;
    dffr camera_module_cache_reg_ram_91__3 (.Q (camera_module_cache_ram_91__3), 
         .QB (\$dummy [1491]), .D (nx9713), .CLK (clk), .R (rst)) ;
    mux21_ni ix9714 (.Y (nx9713), .A0 (camera_module_cache_ram_91__3), .A1 (
             nx35342), .S0 (nx34344)) ;
    aoi22 ix30785 (.Y (nx30784), .A0 (camera_module_cache_ram_123__3), .A1 (
          nx36074), .B0 (camera_module_cache_ram_107__3), .B1 (nx36114)) ;
    dffr camera_module_cache_reg_ram_123__3 (.Q (camera_module_cache_ram_123__3)
         , .QB (\$dummy [1492]), .D (nx9693), .CLK (clk), .R (rst)) ;
    mux21_ni ix9694 (.Y (nx9693), .A0 (camera_module_cache_ram_123__3), .A1 (
             nx35344), .S0 (nx34336)) ;
    dffr camera_module_cache_reg_ram_107__3 (.Q (camera_module_cache_ram_107__3)
         , .QB (\$dummy [1493]), .D (nx9703), .CLK (clk), .R (rst)) ;
    mux21_ni ix9704 (.Y (nx9703), .A0 (camera_module_cache_ram_107__3), .A1 (
             nx35344), .S0 (nx34340)) ;
    nand04 ix12381 (.Y (nx12380), .A0 (nx30793), .A1 (nx30801), .A2 (nx30809), .A3 (
           nx30817)) ;
    aoi22 ix30794 (.Y (nx30793), .A0 (camera_module_cache_ram_139__3), .A1 (
          nx36154), .B0 (camera_module_cache_ram_155__3), .B1 (nx36194)) ;
    dffr camera_module_cache_reg_ram_139__3 (.Q (camera_module_cache_ram_139__3)
         , .QB (\$dummy [1494]), .D (nx9683), .CLK (clk), .R (rst)) ;
    mux21_ni ix9684 (.Y (nx9683), .A0 (camera_module_cache_ram_139__3), .A1 (
             nx35344), .S0 (nx34332)) ;
    dffr camera_module_cache_reg_ram_155__3 (.Q (camera_module_cache_ram_155__3)
         , .QB (\$dummy [1495]), .D (nx9673), .CLK (clk), .R (rst)) ;
    mux21_ni ix9674 (.Y (nx9673), .A0 (camera_module_cache_ram_155__3), .A1 (
             nx35344), .S0 (nx34328)) ;
    aoi22 ix30802 (.Y (nx30801), .A0 (camera_module_cache_ram_187__3), .A1 (
          nx36234), .B0 (camera_module_cache_ram_171__3), .B1 (nx36274)) ;
    dffr camera_module_cache_reg_ram_187__3 (.Q (camera_module_cache_ram_187__3)
         , .QB (\$dummy [1496]), .D (nx9653), .CLK (clk), .R (rst)) ;
    mux21_ni ix9654 (.Y (nx9653), .A0 (camera_module_cache_ram_187__3), .A1 (
             nx35344), .S0 (nx34320)) ;
    dffr camera_module_cache_reg_ram_171__3 (.Q (camera_module_cache_ram_171__3)
         , .QB (\$dummy [1497]), .D (nx9663), .CLK (clk), .R (rst)) ;
    mux21_ni ix9664 (.Y (nx9663), .A0 (camera_module_cache_ram_171__3), .A1 (
             nx35344), .S0 (nx34324)) ;
    aoi22 ix30810 (.Y (nx30809), .A0 (camera_module_cache_ram_203__3), .A1 (
          nx36314), .B0 (camera_module_cache_ram_219__3), .B1 (nx36354)) ;
    dffr camera_module_cache_reg_ram_203__3 (.Q (camera_module_cache_ram_203__3)
         , .QB (\$dummy [1498]), .D (nx9643), .CLK (clk), .R (rst)) ;
    mux21_ni ix9644 (.Y (nx9643), .A0 (camera_module_cache_ram_203__3), .A1 (
             nx35344), .S0 (nx34316)) ;
    dffr camera_module_cache_reg_ram_219__3 (.Q (camera_module_cache_ram_219__3)
         , .QB (\$dummy [1499]), .D (nx9633), .CLK (clk), .R (rst)) ;
    mux21_ni ix9634 (.Y (nx9633), .A0 (camera_module_cache_ram_219__3), .A1 (
             nx35346), .S0 (nx34312)) ;
    aoi22 ix30818 (.Y (nx30817), .A0 (camera_module_cache_ram_235__3), .A1 (
          nx36394), .B0 (camera_module_cache_ram_251__3), .B1 (nx36434)) ;
    dffr camera_module_cache_reg_ram_235__3 (.Q (camera_module_cache_ram_235__3)
         , .QB (\$dummy [1500]), .D (nx9623), .CLK (clk), .R (rst)) ;
    mux21_ni ix9624 (.Y (nx9623), .A0 (camera_module_cache_ram_235__3), .A1 (
             nx35346), .S0 (nx34308)) ;
    dffr camera_module_cache_reg_ram_251__3 (.Q (camera_module_cache_ram_251__3)
         , .QB (\$dummy [1501]), .D (nx9613), .CLK (clk), .R (rst)) ;
    mux21_ni ix9614 (.Y (nx9613), .A0 (camera_module_cache_ram_251__3), .A1 (
             nx35346), .S0 (nx34304)) ;
    nand04 ix12303 (.Y (nx12302), .A0 (nx30826), .A1 (nx30894), .A2 (nx30962), .A3 (
           nx31030)) ;
    oai21 ix30827 (.Y (nx30826), .A0 (nx12292), .A1 (nx12214), .B0 (nx36508)) ;
    nand04 ix12293 (.Y (nx12292), .A0 (nx30829), .A1 (nx30837), .A2 (nx30845), .A3 (
           nx30853)) ;
    aoi22 ix30830 (.Y (nx30829), .A0 (camera_module_cache_ram_12__3), .A1 (
          nx35834), .B0 (camera_module_cache_ram_28__3), .B1 (nx35874)) ;
    dffr camera_module_cache_reg_ram_12__3 (.Q (camera_module_cache_ram_12__3), 
         .QB (\$dummy [1502]), .D (nx9603), .CLK (clk), .R (rst)) ;
    mux21_ni ix9604 (.Y (nx9603), .A0 (nx35346), .A1 (
             camera_module_cache_ram_12__3), .S0 (nx36496)) ;
    dffr camera_module_cache_reg_ram_28__3 (.Q (camera_module_cache_ram_28__3), 
         .QB (\$dummy [1503]), .D (nx9593), .CLK (clk), .R (rst)) ;
    mux21_ni ix9594 (.Y (nx9593), .A0 (nx35346), .A1 (
             camera_module_cache_ram_28__3), .S0 (nx36510)) ;
    aoi22 ix30838 (.Y (nx30837), .A0 (camera_module_cache_ram_44__3), .A1 (
          nx35914), .B0 (camera_module_cache_ram_60__3), .B1 (nx35954)) ;
    dffr camera_module_cache_reg_ram_44__3 (.Q (camera_module_cache_ram_44__3), 
         .QB (\$dummy [1504]), .D (nx9583), .CLK (clk), .R (rst)) ;
    mux21_ni ix9584 (.Y (nx9583), .A0 (nx35346), .A1 (
             camera_module_cache_ram_44__3), .S0 (nx36514)) ;
    dffr camera_module_cache_reg_ram_60__3 (.Q (camera_module_cache_ram_60__3), 
         .QB (\$dummy [1505]), .D (nx9573), .CLK (clk), .R (rst)) ;
    mux21_ni ix9574 (.Y (nx9573), .A0 (nx35346), .A1 (
             camera_module_cache_ram_60__3), .S0 (nx36518)) ;
    aoi22 ix30846 (.Y (nx30845), .A0 (camera_module_cache_ram_76__3), .A1 (
          nx35994), .B0 (camera_module_cache_ram_92__3), .B1 (nx36034)) ;
    dffr camera_module_cache_reg_ram_76__3 (.Q (camera_module_cache_ram_76__3), 
         .QB (\$dummy [1506]), .D (nx9563), .CLK (clk), .R (rst)) ;
    mux21_ni ix9564 (.Y (nx9563), .A0 (nx35348), .A1 (
             camera_module_cache_ram_76__3), .S0 (nx36522)) ;
    dffr camera_module_cache_reg_ram_92__3 (.Q (camera_module_cache_ram_92__3), 
         .QB (\$dummy [1507]), .D (nx9553), .CLK (clk), .R (rst)) ;
    mux21_ni ix9554 (.Y (nx9553), .A0 (nx35348), .A1 (
             camera_module_cache_ram_92__3), .S0 (nx36526)) ;
    aoi22 ix30854 (.Y (nx30853), .A0 (camera_module_cache_ram_124__3), .A1 (
          nx36074), .B0 (camera_module_cache_ram_108__3), .B1 (nx36114)) ;
    dffr camera_module_cache_reg_ram_124__3 (.Q (camera_module_cache_ram_124__3)
         , .QB (\$dummy [1508]), .D (nx9533), .CLK (clk), .R (rst)) ;
    mux21_ni ix9534 (.Y (nx9533), .A0 (nx35348), .A1 (
             camera_module_cache_ram_124__3), .S0 (nx36530)) ;
    dffr camera_module_cache_reg_ram_108__3 (.Q (camera_module_cache_ram_108__3)
         , .QB (\$dummy [1509]), .D (nx9543), .CLK (clk), .R (rst)) ;
    mux21_ni ix9544 (.Y (nx9543), .A0 (nx35348), .A1 (
             camera_module_cache_ram_108__3), .S0 (nx36534)) ;
    nand04 ix12215 (.Y (nx12214), .A0 (nx30862), .A1 (nx30870), .A2 (nx30878), .A3 (
           nx30886)) ;
    aoi22 ix30863 (.Y (nx30862), .A0 (camera_module_cache_ram_140__3), .A1 (
          nx36154), .B0 (camera_module_cache_ram_156__3), .B1 (nx36194)) ;
    dffr camera_module_cache_reg_ram_140__3 (.Q (camera_module_cache_ram_140__3)
         , .QB (\$dummy [1510]), .D (nx9523), .CLK (clk), .R (rst)) ;
    mux21_ni ix9524 (.Y (nx9523), .A0 (nx35348), .A1 (
             camera_module_cache_ram_140__3), .S0 (nx36538)) ;
    dffr camera_module_cache_reg_ram_156__3 (.Q (camera_module_cache_ram_156__3)
         , .QB (\$dummy [1511]), .D (nx9513), .CLK (clk), .R (rst)) ;
    mux21_ni ix9514 (.Y (nx9513), .A0 (nx35348), .A1 (
             camera_module_cache_ram_156__3), .S0 (nx36542)) ;
    aoi22 ix30871 (.Y (nx30870), .A0 (camera_module_cache_ram_188__3), .A1 (
          nx36234), .B0 (camera_module_cache_ram_172__3), .B1 (nx36274)) ;
    dffr camera_module_cache_reg_ram_188__3 (.Q (camera_module_cache_ram_188__3)
         , .QB (\$dummy [1512]), .D (nx9493), .CLK (clk), .R (rst)) ;
    mux21_ni ix9494 (.Y (nx9493), .A0 (nx35348), .A1 (
             camera_module_cache_ram_188__3), .S0 (nx36546)) ;
    dffr camera_module_cache_reg_ram_172__3 (.Q (camera_module_cache_ram_172__3)
         , .QB (\$dummy [1513]), .D (nx9503), .CLK (clk), .R (rst)) ;
    mux21_ni ix9504 (.Y (nx9503), .A0 (nx35350), .A1 (
             camera_module_cache_ram_172__3), .S0 (nx36550)) ;
    aoi22 ix30879 (.Y (nx30878), .A0 (camera_module_cache_ram_204__3), .A1 (
          nx36314), .B0 (camera_module_cache_ram_220__3), .B1 (nx36354)) ;
    dffr camera_module_cache_reg_ram_204__3 (.Q (camera_module_cache_ram_204__3)
         , .QB (\$dummy [1514]), .D (nx9483), .CLK (clk), .R (rst)) ;
    mux21_ni ix9484 (.Y (nx9483), .A0 (nx35350), .A1 (
             camera_module_cache_ram_204__3), .S0 (nx36554)) ;
    dffr camera_module_cache_reg_ram_220__3 (.Q (camera_module_cache_ram_220__3)
         , .QB (\$dummy [1515]), .D (nx9473), .CLK (clk), .R (rst)) ;
    mux21_ni ix9474 (.Y (nx9473), .A0 (nx35350), .A1 (
             camera_module_cache_ram_220__3), .S0 (nx36558)) ;
    aoi22 ix30887 (.Y (nx30886), .A0 (camera_module_cache_ram_236__3), .A1 (
          nx36394), .B0 (camera_module_cache_ram_252__3), .B1 (nx36434)) ;
    dffr camera_module_cache_reg_ram_236__3 (.Q (camera_module_cache_ram_236__3)
         , .QB (\$dummy [1516]), .D (nx9463), .CLK (clk), .R (rst)) ;
    mux21_ni ix9464 (.Y (nx9463), .A0 (nx35350), .A1 (
             camera_module_cache_ram_236__3), .S0 (nx36562)) ;
    dffr camera_module_cache_reg_ram_252__3 (.Q (camera_module_cache_ram_252__3)
         , .QB (\$dummy [1517]), .D (nx9453), .CLK (clk), .R (rst)) ;
    mux21_ni ix9454 (.Y (nx9453), .A0 (nx35350), .A1 (
             camera_module_cache_ram_252__3), .S0 (nx36566)) ;
    oai21 ix30895 (.Y (nx30894), .A0 (nx12130), .A1 (nx12052), .B0 (nx36582)) ;
    nand04 ix12131 (.Y (nx12130), .A0 (nx30897), .A1 (nx30905), .A2 (nx30913), .A3 (
           nx30921)) ;
    aoi22 ix30898 (.Y (nx30897), .A0 (camera_module_cache_ram_13__3), .A1 (
          nx35834), .B0 (camera_module_cache_ram_29__3), .B1 (nx35874)) ;
    dffr camera_module_cache_reg_ram_13__3 (.Q (camera_module_cache_ram_13__3), 
         .QB (\$dummy [1518]), .D (nx9443), .CLK (clk), .R (rst)) ;
    mux21_ni ix9444 (.Y (nx9443), .A0 (nx35350), .A1 (
             camera_module_cache_ram_13__3), .S0 (nx36570)) ;
    dffr camera_module_cache_reg_ram_29__3 (.Q (camera_module_cache_ram_29__3), 
         .QB (\$dummy [1519]), .D (nx9433), .CLK (clk), .R (rst)) ;
    mux21_ni ix9434 (.Y (nx9433), .A0 (nx35350), .A1 (
             camera_module_cache_ram_29__3), .S0 (nx36584)) ;
    aoi22 ix30906 (.Y (nx30905), .A0 (camera_module_cache_ram_45__3), .A1 (
          nx35914), .B0 (camera_module_cache_ram_61__3), .B1 (nx35954)) ;
    dffr camera_module_cache_reg_ram_45__3 (.Q (camera_module_cache_ram_45__3), 
         .QB (\$dummy [1520]), .D (nx9423), .CLK (clk), .R (rst)) ;
    mux21_ni ix9424 (.Y (nx9423), .A0 (nx35352), .A1 (
             camera_module_cache_ram_45__3), .S0 (nx36588)) ;
    dffr camera_module_cache_reg_ram_61__3 (.Q (camera_module_cache_ram_61__3), 
         .QB (\$dummy [1521]), .D (nx9413), .CLK (clk), .R (rst)) ;
    mux21_ni ix9414 (.Y (nx9413), .A0 (nx35352), .A1 (
             camera_module_cache_ram_61__3), .S0 (nx36592)) ;
    aoi22 ix30914 (.Y (nx30913), .A0 (camera_module_cache_ram_77__3), .A1 (
          nx35994), .B0 (camera_module_cache_ram_93__3), .B1 (nx36034)) ;
    dffr camera_module_cache_reg_ram_77__3 (.Q (camera_module_cache_ram_77__3), 
         .QB (\$dummy [1522]), .D (nx9403), .CLK (clk), .R (rst)) ;
    mux21_ni ix9404 (.Y (nx9403), .A0 (nx35352), .A1 (
             camera_module_cache_ram_77__3), .S0 (nx36596)) ;
    dffr camera_module_cache_reg_ram_93__3 (.Q (camera_module_cache_ram_93__3), 
         .QB (\$dummy [1523]), .D (nx9393), .CLK (clk), .R (rst)) ;
    mux21_ni ix9394 (.Y (nx9393), .A0 (nx35352), .A1 (
             camera_module_cache_ram_93__3), .S0 (nx36600)) ;
    aoi22 ix30922 (.Y (nx30921), .A0 (camera_module_cache_ram_125__3), .A1 (
          nx36074), .B0 (camera_module_cache_ram_109__3), .B1 (nx36114)) ;
    dffr camera_module_cache_reg_ram_125__3 (.Q (camera_module_cache_ram_125__3)
         , .QB (\$dummy [1524]), .D (nx9373), .CLK (clk), .R (rst)) ;
    mux21_ni ix9374 (.Y (nx9373), .A0 (nx35352), .A1 (
             camera_module_cache_ram_125__3), .S0 (nx36604)) ;
    dffr camera_module_cache_reg_ram_109__3 (.Q (camera_module_cache_ram_109__3)
         , .QB (\$dummy [1525]), .D (nx9383), .CLK (clk), .R (rst)) ;
    mux21_ni ix9384 (.Y (nx9383), .A0 (nx35352), .A1 (
             camera_module_cache_ram_109__3), .S0 (nx36608)) ;
    nand04 ix12053 (.Y (nx12052), .A0 (nx30930), .A1 (nx30938), .A2 (nx30946), .A3 (
           nx30954)) ;
    aoi22 ix30931 (.Y (nx30930), .A0 (camera_module_cache_ram_141__3), .A1 (
          nx36154), .B0 (camera_module_cache_ram_157__3), .B1 (nx36194)) ;
    dffr camera_module_cache_reg_ram_141__3 (.Q (camera_module_cache_ram_141__3)
         , .QB (\$dummy [1526]), .D (nx9363), .CLK (clk), .R (rst)) ;
    mux21_ni ix9364 (.Y (nx9363), .A0 (nx35352), .A1 (
             camera_module_cache_ram_141__3), .S0 (nx36612)) ;
    dffr camera_module_cache_reg_ram_157__3 (.Q (camera_module_cache_ram_157__3)
         , .QB (\$dummy [1527]), .D (nx9353), .CLK (clk), .R (rst)) ;
    mux21_ni ix9354 (.Y (nx9353), .A0 (nx35354), .A1 (
             camera_module_cache_ram_157__3), .S0 (nx36616)) ;
    aoi22 ix30939 (.Y (nx30938), .A0 (camera_module_cache_ram_189__3), .A1 (
          nx36234), .B0 (camera_module_cache_ram_173__3), .B1 (nx36274)) ;
    dffr camera_module_cache_reg_ram_189__3 (.Q (camera_module_cache_ram_189__3)
         , .QB (\$dummy [1528]), .D (nx9333), .CLK (clk), .R (rst)) ;
    mux21_ni ix9334 (.Y (nx9333), .A0 (nx35354), .A1 (
             camera_module_cache_ram_189__3), .S0 (nx36620)) ;
    dffr camera_module_cache_reg_ram_173__3 (.Q (camera_module_cache_ram_173__3)
         , .QB (\$dummy [1529]), .D (nx9343), .CLK (clk), .R (rst)) ;
    mux21_ni ix9344 (.Y (nx9343), .A0 (nx35354), .A1 (
             camera_module_cache_ram_173__3), .S0 (nx36624)) ;
    aoi22 ix30947 (.Y (nx30946), .A0 (camera_module_cache_ram_205__3), .A1 (
          nx36314), .B0 (camera_module_cache_ram_221__3), .B1 (nx36354)) ;
    dffr camera_module_cache_reg_ram_205__3 (.Q (camera_module_cache_ram_205__3)
         , .QB (\$dummy [1530]), .D (nx9323), .CLK (clk), .R (rst)) ;
    mux21_ni ix9324 (.Y (nx9323), .A0 (nx35354), .A1 (
             camera_module_cache_ram_205__3), .S0 (nx36628)) ;
    dffr camera_module_cache_reg_ram_221__3 (.Q (camera_module_cache_ram_221__3)
         , .QB (\$dummy [1531]), .D (nx9313), .CLK (clk), .R (rst)) ;
    mux21_ni ix9314 (.Y (nx9313), .A0 (nx35354), .A1 (
             camera_module_cache_ram_221__3), .S0 (nx36632)) ;
    aoi22 ix30955 (.Y (nx30954), .A0 (camera_module_cache_ram_237__3), .A1 (
          nx36394), .B0 (camera_module_cache_ram_253__3), .B1 (nx36434)) ;
    dffr camera_module_cache_reg_ram_237__3 (.Q (camera_module_cache_ram_237__3)
         , .QB (\$dummy [1532]), .D (nx9303), .CLK (clk), .R (rst)) ;
    mux21_ni ix9304 (.Y (nx9303), .A0 (nx35354), .A1 (
             camera_module_cache_ram_237__3), .S0 (nx36636)) ;
    dffr camera_module_cache_reg_ram_253__3 (.Q (camera_module_cache_ram_253__3)
         , .QB (\$dummy [1533]), .D (nx9293), .CLK (clk), .R (rst)) ;
    mux21_ni ix9294 (.Y (nx9293), .A0 (nx35354), .A1 (
             camera_module_cache_ram_253__3), .S0 (nx36640)) ;
    oai21 ix30963 (.Y (nx30962), .A0 (nx11966), .A1 (nx11888), .B0 (nx36656)) ;
    nand04 ix11967 (.Y (nx11966), .A0 (nx30965), .A1 (nx30973), .A2 (nx30981), .A3 (
           nx30989)) ;
    aoi22 ix30966 (.Y (nx30965), .A0 (camera_module_cache_ram_14__3), .A1 (
          nx35836), .B0 (camera_module_cache_ram_30__3), .B1 (nx35876)) ;
    dffr camera_module_cache_reg_ram_14__3 (.Q (camera_module_cache_ram_14__3), 
         .QB (\$dummy [1534]), .D (nx9283), .CLK (clk), .R (rst)) ;
    mux21_ni ix9284 (.Y (nx9283), .A0 (nx35356), .A1 (
             camera_module_cache_ram_14__3), .S0 (nx36644)) ;
    dffr camera_module_cache_reg_ram_30__3 (.Q (camera_module_cache_ram_30__3), 
         .QB (\$dummy [1535]), .D (nx9273), .CLK (clk), .R (rst)) ;
    mux21_ni ix9274 (.Y (nx9273), .A0 (nx35356), .A1 (
             camera_module_cache_ram_30__3), .S0 (nx36658)) ;
    aoi22 ix30974 (.Y (nx30973), .A0 (camera_module_cache_ram_46__3), .A1 (
          nx35916), .B0 (camera_module_cache_ram_62__3), .B1 (nx35956)) ;
    dffr camera_module_cache_reg_ram_46__3 (.Q (camera_module_cache_ram_46__3), 
         .QB (\$dummy [1536]), .D (nx9263), .CLK (clk), .R (rst)) ;
    mux21_ni ix9264 (.Y (nx9263), .A0 (nx35356), .A1 (
             camera_module_cache_ram_46__3), .S0 (nx36662)) ;
    dffr camera_module_cache_reg_ram_62__3 (.Q (camera_module_cache_ram_62__3), 
         .QB (\$dummy [1537]), .D (nx9253), .CLK (clk), .R (rst)) ;
    mux21_ni ix9254 (.Y (nx9253), .A0 (nx35356), .A1 (
             camera_module_cache_ram_62__3), .S0 (nx36666)) ;
    aoi22 ix30982 (.Y (nx30981), .A0 (camera_module_cache_ram_78__3), .A1 (
          nx35996), .B0 (camera_module_cache_ram_94__3), .B1 (nx36036)) ;
    dffr camera_module_cache_reg_ram_78__3 (.Q (camera_module_cache_ram_78__3), 
         .QB (\$dummy [1538]), .D (nx9243), .CLK (clk), .R (rst)) ;
    mux21_ni ix9244 (.Y (nx9243), .A0 (nx35356), .A1 (
             camera_module_cache_ram_78__3), .S0 (nx36670)) ;
    dffr camera_module_cache_reg_ram_94__3 (.Q (camera_module_cache_ram_94__3), 
         .QB (\$dummy [1539]), .D (nx9233), .CLK (clk), .R (rst)) ;
    mux21_ni ix9234 (.Y (nx9233), .A0 (nx35356), .A1 (
             camera_module_cache_ram_94__3), .S0 (nx36674)) ;
    aoi22 ix30990 (.Y (nx30989), .A0 (camera_module_cache_ram_126__3), .A1 (
          nx36076), .B0 (camera_module_cache_ram_110__3), .B1 (nx36116)) ;
    dffr camera_module_cache_reg_ram_126__3 (.Q (camera_module_cache_ram_126__3)
         , .QB (\$dummy [1540]), .D (nx9213), .CLK (clk), .R (rst)) ;
    mux21_ni ix9214 (.Y (nx9213), .A0 (nx35356), .A1 (
             camera_module_cache_ram_126__3), .S0 (nx36678)) ;
    dffr camera_module_cache_reg_ram_110__3 (.Q (camera_module_cache_ram_110__3)
         , .QB (\$dummy [1541]), .D (nx9223), .CLK (clk), .R (rst)) ;
    mux21_ni ix9224 (.Y (nx9223), .A0 (nx35358), .A1 (
             camera_module_cache_ram_110__3), .S0 (nx36682)) ;
    nand04 ix11889 (.Y (nx11888), .A0 (nx30998), .A1 (nx31006), .A2 (nx31014), .A3 (
           nx31022)) ;
    aoi22 ix30999 (.Y (nx30998), .A0 (camera_module_cache_ram_142__3), .A1 (
          nx36156), .B0 (camera_module_cache_ram_158__3), .B1 (nx36196)) ;
    dffr camera_module_cache_reg_ram_142__3 (.Q (camera_module_cache_ram_142__3)
         , .QB (\$dummy [1542]), .D (nx9203), .CLK (clk), .R (rst)) ;
    mux21_ni ix9204 (.Y (nx9203), .A0 (nx35358), .A1 (
             camera_module_cache_ram_142__3), .S0 (nx36686)) ;
    dffr camera_module_cache_reg_ram_158__3 (.Q (camera_module_cache_ram_158__3)
         , .QB (\$dummy [1543]), .D (nx9193), .CLK (clk), .R (rst)) ;
    mux21_ni ix9194 (.Y (nx9193), .A0 (nx35358), .A1 (
             camera_module_cache_ram_158__3), .S0 (nx36690)) ;
    aoi22 ix31007 (.Y (nx31006), .A0 (camera_module_cache_ram_190__3), .A1 (
          nx36236), .B0 (camera_module_cache_ram_174__3), .B1 (nx36276)) ;
    dffr camera_module_cache_reg_ram_190__3 (.Q (camera_module_cache_ram_190__3)
         , .QB (\$dummy [1544]), .D (nx9173), .CLK (clk), .R (rst)) ;
    mux21_ni ix9174 (.Y (nx9173), .A0 (nx35358), .A1 (
             camera_module_cache_ram_190__3), .S0 (nx36694)) ;
    dffr camera_module_cache_reg_ram_174__3 (.Q (camera_module_cache_ram_174__3)
         , .QB (\$dummy [1545]), .D (nx9183), .CLK (clk), .R (rst)) ;
    mux21_ni ix9184 (.Y (nx9183), .A0 (nx35358), .A1 (
             camera_module_cache_ram_174__3), .S0 (nx36698)) ;
    aoi22 ix31015 (.Y (nx31014), .A0 (camera_module_cache_ram_206__3), .A1 (
          nx36316), .B0 (camera_module_cache_ram_222__3), .B1 (nx36356)) ;
    dffr camera_module_cache_reg_ram_206__3 (.Q (camera_module_cache_ram_206__3)
         , .QB (\$dummy [1546]), .D (nx9163), .CLK (clk), .R (rst)) ;
    mux21_ni ix9164 (.Y (nx9163), .A0 (nx35358), .A1 (
             camera_module_cache_ram_206__3), .S0 (nx36702)) ;
    dffr camera_module_cache_reg_ram_222__3 (.Q (camera_module_cache_ram_222__3)
         , .QB (\$dummy [1547]), .D (nx9153), .CLK (clk), .R (rst)) ;
    mux21_ni ix9154 (.Y (nx9153), .A0 (nx35358), .A1 (
             camera_module_cache_ram_222__3), .S0 (nx36706)) ;
    aoi22 ix31023 (.Y (nx31022), .A0 (camera_module_cache_ram_238__3), .A1 (
          nx36396), .B0 (camera_module_cache_ram_254__3), .B1 (nx36436)) ;
    dffr camera_module_cache_reg_ram_238__3 (.Q (camera_module_cache_ram_238__3)
         , .QB (\$dummy [1548]), .D (nx9143), .CLK (clk), .R (rst)) ;
    mux21_ni ix9144 (.Y (nx9143), .A0 (nx35360), .A1 (
             camera_module_cache_ram_238__3), .S0 (nx36710)) ;
    dffr camera_module_cache_reg_ram_254__3 (.Q (camera_module_cache_ram_254__3)
         , .QB (\$dummy [1549]), .D (nx9133), .CLK (clk), .R (rst)) ;
    mux21_ni ix9134 (.Y (nx9133), .A0 (nx35360), .A1 (
             camera_module_cache_ram_254__3), .S0 (nx36714)) ;
    oai21 ix31031 (.Y (nx31030), .A0 (nx11804), .A1 (nx11726), .B0 (nx36730)) ;
    nand04 ix11805 (.Y (nx11804), .A0 (nx31033), .A1 (nx31041), .A2 (nx31049), .A3 (
           nx31057)) ;
    aoi22 ix31034 (.Y (nx31033), .A0 (camera_module_cache_ram_15__3), .A1 (
          nx35836), .B0 (camera_module_cache_ram_31__3), .B1 (nx35876)) ;
    dffr camera_module_cache_reg_ram_15__3 (.Q (camera_module_cache_ram_15__3), 
         .QB (\$dummy [1550]), .D (nx9123), .CLK (clk), .R (rst)) ;
    mux21_ni ix9124 (.Y (nx9123), .A0 (nx35360), .A1 (
             camera_module_cache_ram_15__3), .S0 (nx36718)) ;
    dffr camera_module_cache_reg_ram_31__3 (.Q (camera_module_cache_ram_31__3), 
         .QB (\$dummy [1551]), .D (nx9113), .CLK (clk), .R (rst)) ;
    mux21_ni ix9114 (.Y (nx9113), .A0 (nx35360), .A1 (
             camera_module_cache_ram_31__3), .S0 (nx36732)) ;
    aoi22 ix31042 (.Y (nx31041), .A0 (camera_module_cache_ram_47__3), .A1 (
          nx35916), .B0 (camera_module_cache_ram_63__3), .B1 (nx35956)) ;
    dffr camera_module_cache_reg_ram_47__3 (.Q (camera_module_cache_ram_47__3), 
         .QB (\$dummy [1552]), .D (nx9103), .CLK (clk), .R (rst)) ;
    mux21_ni ix9104 (.Y (nx9103), .A0 (nx35360), .A1 (
             camera_module_cache_ram_47__3), .S0 (nx36736)) ;
    dffr camera_module_cache_reg_ram_63__3 (.Q (camera_module_cache_ram_63__3), 
         .QB (\$dummy [1553]), .D (nx9093), .CLK (clk), .R (rst)) ;
    mux21_ni ix9094 (.Y (nx9093), .A0 (nx35360), .A1 (
             camera_module_cache_ram_63__3), .S0 (nx36740)) ;
    aoi22 ix31050 (.Y (nx31049), .A0 (camera_module_cache_ram_79__3), .A1 (
          nx35996), .B0 (camera_module_cache_ram_95__3), .B1 (nx36036)) ;
    dffr camera_module_cache_reg_ram_79__3 (.Q (camera_module_cache_ram_79__3), 
         .QB (\$dummy [1554]), .D (nx9083), .CLK (clk), .R (rst)) ;
    mux21_ni ix9084 (.Y (nx9083), .A0 (nx35360), .A1 (
             camera_module_cache_ram_79__3), .S0 (nx36744)) ;
    dffr camera_module_cache_reg_ram_95__3 (.Q (camera_module_cache_ram_95__3), 
         .QB (\$dummy [1555]), .D (nx9073), .CLK (clk), .R (rst)) ;
    mux21_ni ix9074 (.Y (nx9073), .A0 (nx35362), .A1 (
             camera_module_cache_ram_95__3), .S0 (nx36748)) ;
    aoi22 ix31058 (.Y (nx31057), .A0 (camera_module_cache_ram_127__3), .A1 (
          nx36076), .B0 (camera_module_cache_ram_111__3), .B1 (nx36116)) ;
    dffr camera_module_cache_reg_ram_127__3 (.Q (camera_module_cache_ram_127__3)
         , .QB (\$dummy [1556]), .D (nx9053), .CLK (clk), .R (rst)) ;
    mux21_ni ix9054 (.Y (nx9053), .A0 (nx35362), .A1 (
             camera_module_cache_ram_127__3), .S0 (nx36752)) ;
    dffr camera_module_cache_reg_ram_111__3 (.Q (camera_module_cache_ram_111__3)
         , .QB (\$dummy [1557]), .D (nx9063), .CLK (clk), .R (rst)) ;
    mux21_ni ix9064 (.Y (nx9063), .A0 (nx35362), .A1 (
             camera_module_cache_ram_111__3), .S0 (nx36756)) ;
    nand04 ix11727 (.Y (nx11726), .A0 (nx31066), .A1 (nx31074), .A2 (nx31082), .A3 (
           nx31090)) ;
    aoi22 ix31067 (.Y (nx31066), .A0 (camera_module_cache_ram_143__3), .A1 (
          nx36156), .B0 (camera_module_cache_ram_159__3), .B1 (nx36196)) ;
    dffr camera_module_cache_reg_ram_143__3 (.Q (camera_module_cache_ram_143__3)
         , .QB (\$dummy [1558]), .D (nx9043), .CLK (clk), .R (rst)) ;
    mux21_ni ix9044 (.Y (nx9043), .A0 (nx35362), .A1 (
             camera_module_cache_ram_143__3), .S0 (nx36760)) ;
    dffr camera_module_cache_reg_ram_159__3 (.Q (camera_module_cache_ram_159__3)
         , .QB (\$dummy [1559]), .D (nx9033), .CLK (clk), .R (rst)) ;
    mux21_ni ix9034 (.Y (nx9033), .A0 (nx35362), .A1 (
             camera_module_cache_ram_159__3), .S0 (nx36764)) ;
    aoi22 ix31075 (.Y (nx31074), .A0 (camera_module_cache_ram_191__3), .A1 (
          nx36236), .B0 (camera_module_cache_ram_175__3), .B1 (nx36276)) ;
    dffr camera_module_cache_reg_ram_191__3 (.Q (camera_module_cache_ram_191__3)
         , .QB (\$dummy [1560]), .D (nx9013), .CLK (clk), .R (rst)) ;
    mux21_ni ix9014 (.Y (nx9013), .A0 (nx35362), .A1 (
             camera_module_cache_ram_191__3), .S0 (nx36768)) ;
    dffr camera_module_cache_reg_ram_175__3 (.Q (camera_module_cache_ram_175__3)
         , .QB (\$dummy [1561]), .D (nx9023), .CLK (clk), .R (rst)) ;
    mux21_ni ix9024 (.Y (nx9023), .A0 (nx35362), .A1 (
             camera_module_cache_ram_175__3), .S0 (nx36772)) ;
    aoi22 ix31083 (.Y (nx31082), .A0 (camera_module_cache_ram_207__3), .A1 (
          nx36316), .B0 (camera_module_cache_ram_223__3), .B1 (nx36356)) ;
    dffr camera_module_cache_reg_ram_207__3 (.Q (camera_module_cache_ram_207__3)
         , .QB (\$dummy [1562]), .D (nx9003), .CLK (clk), .R (rst)) ;
    mux21_ni ix9004 (.Y (nx9003), .A0 (nx35364), .A1 (
             camera_module_cache_ram_207__3), .S0 (nx36776)) ;
    dffr camera_module_cache_reg_ram_223__3 (.Q (camera_module_cache_ram_223__3)
         , .QB (\$dummy [1563]), .D (nx8993), .CLK (clk), .R (rst)) ;
    mux21_ni ix8994 (.Y (nx8993), .A0 (nx35364), .A1 (
             camera_module_cache_ram_223__3), .S0 (nx36780)) ;
    aoi22 ix31091 (.Y (nx31090), .A0 (camera_module_cache_ram_239__3), .A1 (
          nx36396), .B0 (camera_module_cache_ram_255__3), .B1 (nx36436)) ;
    dffr camera_module_cache_reg_ram_239__3 (.Q (camera_module_cache_ram_239__3)
         , .QB (\$dummy [1564]), .D (nx8983), .CLK (clk), .R (rst)) ;
    mux21_ni ix8984 (.Y (nx8983), .A0 (nx35364), .A1 (
             camera_module_cache_ram_239__3), .S0 (nx36784)) ;
    dffr camera_module_cache_reg_ram_255__3 (.Q (camera_module_cache_ram_255__3)
         , .QB (\$dummy [1565]), .D (nx8973), .CLK (clk), .R (rst)) ;
    mux21_ni ix8974 (.Y (nx8973), .A0 (nx35364), .A1 (
             camera_module_cache_ram_255__3), .S0 (nx36788)) ;
    dff camera_module_algo_module_pixel_reg_reg_q_5 (.Q (
        camera_module_algo_module_pixel_value_5), .QB (nx32240), .D (nx16673), .CLK (
        clk)) ;
    mux21_ni ix16674 (.Y (nx16673), .A0 (nx19834), .A1 (
             camera_module_algo_module_pixel_value_5), .S0 (nx22665)) ;
    mux21_ni ix31107 (.Y (nx31106), .A0 (nx31108), .A1 (nx35676), .S0 (nx36792)
             ) ;
    nor04 ix31109 (.Y (nx31108), .A0 (nx19814), .A1 (nx19160), .A2 (nx18504), .A3 (
          nx17850)) ;
    nand04 ix19815 (.Y (nx19814), .A0 (nx31111), .A1 (nx31217), .A2 (nx31285), .A3 (
           nx31353)) ;
    oai21 ix31112 (.Y (nx31111), .A0 (nx19804), .A1 (nx19726), .B0 (nx36448)) ;
    nand04 ix19805 (.Y (nx19804), .A0 (nx31114), .A1 (nx31160), .A2 (nx31168), .A3 (
           nx31176)) ;
    aoi22 ix31115 (.Y (nx31114), .A0 (camera_module_cache_ram_0__5), .A1 (
          nx35836), .B0 (camera_module_cache_ram_16__5), .B1 (nx35876)) ;
    dffr camera_module_cache_reg_ram_0__5 (.Q (camera_module_cache_ram_0__5), .QB (
         \$dummy [1566]), .D (nx16663), .CLK (clk), .R (rst)) ;
    mux21_ni ix16664 (.Y (nx16663), .A0 (camera_module_cache_ram_0__5), .A1 (
             nx35444), .S0 (nx35134)) ;
    oai221 ix17197 (.Y (nx17196), .A0 (nx34076), .A1 (nx31119), .B0 (nx31135), .B1 (
           nx35714), .C0 (nx31138)) ;
    tri01 nvm_module_tri_dataout_125 (.Y (nvm_data_125), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_117 (.Y (nvm_data_117), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_109 (.Y (nvm_data_109), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_101 (.Y (nvm_data_101), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_93 (.Y (nvm_data_93), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_85 (.Y (nvm_data_85), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_77 (.Y (nvm_data_77), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_69 (.Y (nvm_data_69), .A (nx22549), .E (
          nvm_module_GND0)) ;
    inv01 ix31136 (.Y (nx31135), .A (nvm_data_5)) ;
    tri01 nvm_module_tri_dataout_5 (.Y (nvm_data_5), .A (nx22549), .E (
          nvm_module_GND0)) ;
    nand02 ix31139 (.Y (nx31138), .A0 (nx34076), .A1 (nx17130)) ;
    tri01 nvm_module_tri_dataout_61 (.Y (nvm_data_61), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_53 (.Y (nvm_data_53), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_45 (.Y (nvm_data_45), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_37 (.Y (nvm_data_37), .A (nx22549), .E (
          nvm_module_GND0)) ;
    oai22 ix17099 (.Y (nx17098), .A0 (nx34108), .A1 (nx31149), .B0 (nx34094), .B1 (
          nx31153)) ;
    tri01 nvm_module_tri_dataout_29 (.Y (nvm_data_29), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_21 (.Y (nvm_data_21), .A (nx22549), .E (
          nvm_module_GND0)) ;
    nand02 ix31154 (.Y (nx31153), .A0 (nvm_data_13), .A1 (nx34108)) ;
    tri01 nvm_module_tri_dataout_13 (.Y (nvm_data_13), .A (nx22549), .E (
          nvm_module_GND0)) ;
    dffr camera_module_cache_reg_ram_16__5 (.Q (camera_module_cache_ram_16__5), 
         .QB (\$dummy [1567]), .D (nx16653), .CLK (clk), .R (rst)) ;
    mux21_ni ix16654 (.Y (nx16653), .A0 (camera_module_cache_ram_16__5), .A1 (
             nx35444), .S0 (nx35130)) ;
    aoi22 ix31161 (.Y (nx31160), .A0 (camera_module_cache_ram_32__5), .A1 (
          nx35916), .B0 (camera_module_cache_ram_48__5), .B1 (nx35956)) ;
    dffr camera_module_cache_reg_ram_32__5 (.Q (camera_module_cache_ram_32__5), 
         .QB (\$dummy [1568]), .D (nx16643), .CLK (clk), .R (rst)) ;
    mux21_ni ix16644 (.Y (nx16643), .A0 (camera_module_cache_ram_32__5), .A1 (
             nx35444), .S0 (nx35126)) ;
    dffr camera_module_cache_reg_ram_48__5 (.Q (camera_module_cache_ram_48__5), 
         .QB (\$dummy [1569]), .D (nx16633), .CLK (clk), .R (rst)) ;
    mux21_ni ix16634 (.Y (nx16633), .A0 (camera_module_cache_ram_48__5), .A1 (
             nx35444), .S0 (nx35122)) ;
    aoi22 ix31169 (.Y (nx31168), .A0 (camera_module_cache_ram_64__5), .A1 (
          nx35996), .B0 (camera_module_cache_ram_80__5), .B1 (nx36036)) ;
    dffr camera_module_cache_reg_ram_64__5 (.Q (camera_module_cache_ram_64__5), 
         .QB (\$dummy [1570]), .D (nx16623), .CLK (clk), .R (rst)) ;
    mux21_ni ix16624 (.Y (nx16623), .A0 (camera_module_cache_ram_64__5), .A1 (
             nx35444), .S0 (nx35118)) ;
    dffr camera_module_cache_reg_ram_80__5 (.Q (camera_module_cache_ram_80__5), 
         .QB (\$dummy [1571]), .D (nx16613), .CLK (clk), .R (rst)) ;
    mux21_ni ix16614 (.Y (nx16613), .A0 (camera_module_cache_ram_80__5), .A1 (
             nx35444), .S0 (nx35114)) ;
    aoi22 ix31177 (.Y (nx31176), .A0 (camera_module_cache_ram_112__5), .A1 (
          nx36076), .B0 (camera_module_cache_ram_96__5), .B1 (nx36116)) ;
    dffr camera_module_cache_reg_ram_112__5 (.Q (camera_module_cache_ram_112__5)
         , .QB (\$dummy [1572]), .D (nx16593), .CLK (clk), .R (rst)) ;
    mux21_ni ix16594 (.Y (nx16593), .A0 (camera_module_cache_ram_112__5), .A1 (
             nx35444), .S0 (nx35106)) ;
    dffr camera_module_cache_reg_ram_96__5 (.Q (camera_module_cache_ram_96__5), 
         .QB (\$dummy [1573]), .D (nx16603), .CLK (clk), .R (rst)) ;
    mux21_ni ix16604 (.Y (nx16603), .A0 (camera_module_cache_ram_96__5), .A1 (
             nx35446), .S0 (nx35110)) ;
    nand04 ix19727 (.Y (nx19726), .A0 (nx31185), .A1 (nx31193), .A2 (nx31201), .A3 (
           nx31209)) ;
    aoi22 ix31186 (.Y (nx31185), .A0 (camera_module_cache_ram_128__5), .A1 (
          nx36156), .B0 (camera_module_cache_ram_144__5), .B1 (nx36196)) ;
    dffr camera_module_cache_reg_ram_128__5 (.Q (camera_module_cache_ram_128__5)
         , .QB (\$dummy [1574]), .D (nx16583), .CLK (clk), .R (rst)) ;
    mux21_ni ix16584 (.Y (nx16583), .A0 (camera_module_cache_ram_128__5), .A1 (
             nx35446), .S0 (nx35102)) ;
    dffr camera_module_cache_reg_ram_144__5 (.Q (camera_module_cache_ram_144__5)
         , .QB (\$dummy [1575]), .D (nx16573), .CLK (clk), .R (rst)) ;
    mux21_ni ix16574 (.Y (nx16573), .A0 (camera_module_cache_ram_144__5), .A1 (
             nx35446), .S0 (nx35098)) ;
    aoi22 ix31194 (.Y (nx31193), .A0 (camera_module_cache_ram_176__5), .A1 (
          nx36236), .B0 (camera_module_cache_ram_160__5), .B1 (nx36276)) ;
    dffr camera_module_cache_reg_ram_176__5 (.Q (camera_module_cache_ram_176__5)
         , .QB (\$dummy [1576]), .D (nx16553), .CLK (clk), .R (rst)) ;
    mux21_ni ix16554 (.Y (nx16553), .A0 (camera_module_cache_ram_176__5), .A1 (
             nx35446), .S0 (nx35090)) ;
    dffr camera_module_cache_reg_ram_160__5 (.Q (camera_module_cache_ram_160__5)
         , .QB (\$dummy [1577]), .D (nx16563), .CLK (clk), .R (rst)) ;
    mux21_ni ix16564 (.Y (nx16563), .A0 (camera_module_cache_ram_160__5), .A1 (
             nx35446), .S0 (nx35094)) ;
    aoi22 ix31202 (.Y (nx31201), .A0 (camera_module_cache_ram_192__5), .A1 (
          nx36316), .B0 (camera_module_cache_ram_208__5), .B1 (nx36356)) ;
    dffr camera_module_cache_reg_ram_192__5 (.Q (camera_module_cache_ram_192__5)
         , .QB (\$dummy [1578]), .D (nx16543), .CLK (clk), .R (rst)) ;
    mux21_ni ix16544 (.Y (nx16543), .A0 (camera_module_cache_ram_192__5), .A1 (
             nx35446), .S0 (nx35086)) ;
    dffr camera_module_cache_reg_ram_208__5 (.Q (camera_module_cache_ram_208__5)
         , .QB (\$dummy [1579]), .D (nx16533), .CLK (clk), .R (rst)) ;
    mux21_ni ix16534 (.Y (nx16533), .A0 (camera_module_cache_ram_208__5), .A1 (
             nx35446), .S0 (nx35082)) ;
    aoi22 ix31210 (.Y (nx31209), .A0 (camera_module_cache_ram_224__5), .A1 (
          nx36396), .B0 (camera_module_cache_ram_240__5), .B1 (nx36436)) ;
    dffr camera_module_cache_reg_ram_224__5 (.Q (camera_module_cache_ram_224__5)
         , .QB (\$dummy [1580]), .D (nx16523), .CLK (clk), .R (rst)) ;
    mux21_ni ix16524 (.Y (nx16523), .A0 (camera_module_cache_ram_224__5), .A1 (
             nx35448), .S0 (nx35078)) ;
    dffr camera_module_cache_reg_ram_240__5 (.Q (camera_module_cache_ram_240__5)
         , .QB (\$dummy [1581]), .D (nx16513), .CLK (clk), .R (rst)) ;
    mux21_ni ix16514 (.Y (nx16513), .A0 (camera_module_cache_ram_240__5), .A1 (
             nx35448), .S0 (nx35074)) ;
    oai21 ix31218 (.Y (nx31217), .A0 (nx19642), .A1 (nx19564), .B0 (nx36452)) ;
    nand04 ix19643 (.Y (nx19642), .A0 (nx31220), .A1 (nx31228), .A2 (nx31236), .A3 (
           nx31244)) ;
    aoi22 ix31221 (.Y (nx31220), .A0 (camera_module_cache_ram_1__5), .A1 (
          nx35836), .B0 (camera_module_cache_ram_17__5), .B1 (nx35876)) ;
    dffr camera_module_cache_reg_ram_1__5 (.Q (camera_module_cache_ram_1__5), .QB (
         \$dummy [1582]), .D (nx16503), .CLK (clk), .R (rst)) ;
    mux21_ni ix16504 (.Y (nx16503), .A0 (camera_module_cache_ram_1__5), .A1 (
             nx35448), .S0 (nx35064)) ;
    dffr camera_module_cache_reg_ram_17__5 (.Q (camera_module_cache_ram_17__5), 
         .QB (\$dummy [1583]), .D (nx16493), .CLK (clk), .R (rst)) ;
    mux21_ni ix16494 (.Y (nx16493), .A0 (camera_module_cache_ram_17__5), .A1 (
             nx35448), .S0 (nx35060)) ;
    aoi22 ix31229 (.Y (nx31228), .A0 (camera_module_cache_ram_33__5), .A1 (
          nx35916), .B0 (camera_module_cache_ram_49__5), .B1 (nx35956)) ;
    dffr camera_module_cache_reg_ram_33__5 (.Q (camera_module_cache_ram_33__5), 
         .QB (\$dummy [1584]), .D (nx16483), .CLK (clk), .R (rst)) ;
    mux21_ni ix16484 (.Y (nx16483), .A0 (camera_module_cache_ram_33__5), .A1 (
             nx35448), .S0 (nx35056)) ;
    dffr camera_module_cache_reg_ram_49__5 (.Q (camera_module_cache_ram_49__5), 
         .QB (\$dummy [1585]), .D (nx16473), .CLK (clk), .R (rst)) ;
    mux21_ni ix16474 (.Y (nx16473), .A0 (camera_module_cache_ram_49__5), .A1 (
             nx35448), .S0 (nx35052)) ;
    aoi22 ix31237 (.Y (nx31236), .A0 (camera_module_cache_ram_65__5), .A1 (
          nx35996), .B0 (camera_module_cache_ram_81__5), .B1 (nx36036)) ;
    dffr camera_module_cache_reg_ram_65__5 (.Q (camera_module_cache_ram_65__5), 
         .QB (\$dummy [1586]), .D (nx16463), .CLK (clk), .R (rst)) ;
    mux21_ni ix16464 (.Y (nx16463), .A0 (camera_module_cache_ram_65__5), .A1 (
             nx35448), .S0 (nx35048)) ;
    dffr camera_module_cache_reg_ram_81__5 (.Q (camera_module_cache_ram_81__5), 
         .QB (\$dummy [1587]), .D (nx16453), .CLK (clk), .R (rst)) ;
    mux21_ni ix16454 (.Y (nx16453), .A0 (camera_module_cache_ram_81__5), .A1 (
             nx35450), .S0 (nx35044)) ;
    aoi22 ix31245 (.Y (nx31244), .A0 (camera_module_cache_ram_113__5), .A1 (
          nx36076), .B0 (camera_module_cache_ram_97__5), .B1 (nx36116)) ;
    dffr camera_module_cache_reg_ram_113__5 (.Q (camera_module_cache_ram_113__5)
         , .QB (\$dummy [1588]), .D (nx16433), .CLK (clk), .R (rst)) ;
    mux21_ni ix16434 (.Y (nx16433), .A0 (camera_module_cache_ram_113__5), .A1 (
             nx35450), .S0 (nx35036)) ;
    dffr camera_module_cache_reg_ram_97__5 (.Q (camera_module_cache_ram_97__5), 
         .QB (\$dummy [1589]), .D (nx16443), .CLK (clk), .R (rst)) ;
    mux21_ni ix16444 (.Y (nx16443), .A0 (camera_module_cache_ram_97__5), .A1 (
             nx35450), .S0 (nx35040)) ;
    nand04 ix19565 (.Y (nx19564), .A0 (nx31253), .A1 (nx31261), .A2 (nx31269), .A3 (
           nx31277)) ;
    aoi22 ix31254 (.Y (nx31253), .A0 (camera_module_cache_ram_129__5), .A1 (
          nx36156), .B0 (camera_module_cache_ram_145__5), .B1 (nx36196)) ;
    dffr camera_module_cache_reg_ram_129__5 (.Q (camera_module_cache_ram_129__5)
         , .QB (\$dummy [1590]), .D (nx16423), .CLK (clk), .R (rst)) ;
    mux21_ni ix16424 (.Y (nx16423), .A0 (camera_module_cache_ram_129__5), .A1 (
             nx35450), .S0 (nx35032)) ;
    dffr camera_module_cache_reg_ram_145__5 (.Q (camera_module_cache_ram_145__5)
         , .QB (\$dummy [1591]), .D (nx16413), .CLK (clk), .R (rst)) ;
    mux21_ni ix16414 (.Y (nx16413), .A0 (camera_module_cache_ram_145__5), .A1 (
             nx35450), .S0 (nx35028)) ;
    aoi22 ix31262 (.Y (nx31261), .A0 (camera_module_cache_ram_177__5), .A1 (
          nx36236), .B0 (camera_module_cache_ram_161__5), .B1 (nx36276)) ;
    dffr camera_module_cache_reg_ram_177__5 (.Q (camera_module_cache_ram_177__5)
         , .QB (\$dummy [1592]), .D (nx16393), .CLK (clk), .R (rst)) ;
    mux21_ni ix16394 (.Y (nx16393), .A0 (camera_module_cache_ram_177__5), .A1 (
             nx35450), .S0 (nx35020)) ;
    dffr camera_module_cache_reg_ram_161__5 (.Q (camera_module_cache_ram_161__5)
         , .QB (\$dummy [1593]), .D (nx16403), .CLK (clk), .R (rst)) ;
    mux21_ni ix16404 (.Y (nx16403), .A0 (camera_module_cache_ram_161__5), .A1 (
             nx35450), .S0 (nx35024)) ;
    aoi22 ix31270 (.Y (nx31269), .A0 (camera_module_cache_ram_193__5), .A1 (
          nx36316), .B0 (camera_module_cache_ram_209__5), .B1 (nx36356)) ;
    dffr camera_module_cache_reg_ram_193__5 (.Q (camera_module_cache_ram_193__5)
         , .QB (\$dummy [1594]), .D (nx16383), .CLK (clk), .R (rst)) ;
    mux21_ni ix16384 (.Y (nx16383), .A0 (camera_module_cache_ram_193__5), .A1 (
             nx35452), .S0 (nx35016)) ;
    dffr camera_module_cache_reg_ram_209__5 (.Q (camera_module_cache_ram_209__5)
         , .QB (\$dummy [1595]), .D (nx16373), .CLK (clk), .R (rst)) ;
    mux21_ni ix16374 (.Y (nx16373), .A0 (camera_module_cache_ram_209__5), .A1 (
             nx35452), .S0 (nx35012)) ;
    aoi22 ix31278 (.Y (nx31277), .A0 (camera_module_cache_ram_225__5), .A1 (
          nx36396), .B0 (camera_module_cache_ram_241__5), .B1 (nx36436)) ;
    dffr camera_module_cache_reg_ram_225__5 (.Q (camera_module_cache_ram_225__5)
         , .QB (\$dummy [1596]), .D (nx16363), .CLK (clk), .R (rst)) ;
    mux21_ni ix16364 (.Y (nx16363), .A0 (camera_module_cache_ram_225__5), .A1 (
             nx35452), .S0 (nx35008)) ;
    dffr camera_module_cache_reg_ram_241__5 (.Q (camera_module_cache_ram_241__5)
         , .QB (\$dummy [1597]), .D (nx16353), .CLK (clk), .R (rst)) ;
    mux21_ni ix16354 (.Y (nx16353), .A0 (camera_module_cache_ram_241__5), .A1 (
             nx35452), .S0 (nx35004)) ;
    oai21 ix31286 (.Y (nx31285), .A0 (nx19478), .A1 (nx19400), .B0 (nx36456)) ;
    nand04 ix19479 (.Y (nx19478), .A0 (nx31288), .A1 (nx31296), .A2 (nx31304), .A3 (
           nx31312)) ;
    aoi22 ix31289 (.Y (nx31288), .A0 (camera_module_cache_ram_2__5), .A1 (
          nx35836), .B0 (camera_module_cache_ram_18__5), .B1 (nx35876)) ;
    dffr camera_module_cache_reg_ram_2__5 (.Q (camera_module_cache_ram_2__5), .QB (
         \$dummy [1598]), .D (nx16343), .CLK (clk), .R (rst)) ;
    mux21_ni ix16344 (.Y (nx16343), .A0 (camera_module_cache_ram_2__5), .A1 (
             nx35452), .S0 (nx34994)) ;
    dffr camera_module_cache_reg_ram_18__5 (.Q (camera_module_cache_ram_18__5), 
         .QB (\$dummy [1599]), .D (nx16333), .CLK (clk), .R (rst)) ;
    mux21_ni ix16334 (.Y (nx16333), .A0 (camera_module_cache_ram_18__5), .A1 (
             nx35452), .S0 (nx34990)) ;
    aoi22 ix31297 (.Y (nx31296), .A0 (camera_module_cache_ram_34__5), .A1 (
          nx35916), .B0 (camera_module_cache_ram_50__5), .B1 (nx35956)) ;
    dffr camera_module_cache_reg_ram_34__5 (.Q (camera_module_cache_ram_34__5), 
         .QB (\$dummy [1600]), .D (nx16323), .CLK (clk), .R (rst)) ;
    mux21_ni ix16324 (.Y (nx16323), .A0 (camera_module_cache_ram_34__5), .A1 (
             nx35452), .S0 (nx34986)) ;
    dffr camera_module_cache_reg_ram_50__5 (.Q (camera_module_cache_ram_50__5), 
         .QB (\$dummy [1601]), .D (nx16313), .CLK (clk), .R (rst)) ;
    mux21_ni ix16314 (.Y (nx16313), .A0 (camera_module_cache_ram_50__5), .A1 (
             nx35454), .S0 (nx34982)) ;
    aoi22 ix31305 (.Y (nx31304), .A0 (camera_module_cache_ram_66__5), .A1 (
          nx35996), .B0 (camera_module_cache_ram_82__5), .B1 (nx36036)) ;
    dffr camera_module_cache_reg_ram_66__5 (.Q (camera_module_cache_ram_66__5), 
         .QB (\$dummy [1602]), .D (nx16303), .CLK (clk), .R (rst)) ;
    mux21_ni ix16304 (.Y (nx16303), .A0 (camera_module_cache_ram_66__5), .A1 (
             nx35454), .S0 (nx34978)) ;
    dffr camera_module_cache_reg_ram_82__5 (.Q (camera_module_cache_ram_82__5), 
         .QB (\$dummy [1603]), .D (nx16293), .CLK (clk), .R (rst)) ;
    mux21_ni ix16294 (.Y (nx16293), .A0 (camera_module_cache_ram_82__5), .A1 (
             nx35454), .S0 (nx34974)) ;
    aoi22 ix31313 (.Y (nx31312), .A0 (camera_module_cache_ram_114__5), .A1 (
          nx36076), .B0 (camera_module_cache_ram_98__5), .B1 (nx36116)) ;
    dffr camera_module_cache_reg_ram_114__5 (.Q (camera_module_cache_ram_114__5)
         , .QB (\$dummy [1604]), .D (nx16273), .CLK (clk), .R (rst)) ;
    mux21_ni ix16274 (.Y (nx16273), .A0 (camera_module_cache_ram_114__5), .A1 (
             nx35454), .S0 (nx34966)) ;
    dffr camera_module_cache_reg_ram_98__5 (.Q (camera_module_cache_ram_98__5), 
         .QB (\$dummy [1605]), .D (nx16283), .CLK (clk), .R (rst)) ;
    mux21_ni ix16284 (.Y (nx16283), .A0 (camera_module_cache_ram_98__5), .A1 (
             nx35454), .S0 (nx34970)) ;
    nand04 ix19401 (.Y (nx19400), .A0 (nx31321), .A1 (nx31329), .A2 (nx31337), .A3 (
           nx31345)) ;
    aoi22 ix31322 (.Y (nx31321), .A0 (camera_module_cache_ram_130__5), .A1 (
          nx36156), .B0 (camera_module_cache_ram_146__5), .B1 (nx36196)) ;
    dffr camera_module_cache_reg_ram_130__5 (.Q (camera_module_cache_ram_130__5)
         , .QB (\$dummy [1606]), .D (nx16263), .CLK (clk), .R (rst)) ;
    mux21_ni ix16264 (.Y (nx16263), .A0 (camera_module_cache_ram_130__5), .A1 (
             nx35454), .S0 (nx34962)) ;
    dffr camera_module_cache_reg_ram_146__5 (.Q (camera_module_cache_ram_146__5)
         , .QB (\$dummy [1607]), .D (nx16253), .CLK (clk), .R (rst)) ;
    mux21_ni ix16254 (.Y (nx16253), .A0 (camera_module_cache_ram_146__5), .A1 (
             nx35454), .S0 (nx34958)) ;
    aoi22 ix31330 (.Y (nx31329), .A0 (camera_module_cache_ram_178__5), .A1 (
          nx36236), .B0 (camera_module_cache_ram_162__5), .B1 (nx36276)) ;
    dffr camera_module_cache_reg_ram_178__5 (.Q (camera_module_cache_ram_178__5)
         , .QB (\$dummy [1608]), .D (nx16233), .CLK (clk), .R (rst)) ;
    mux21_ni ix16234 (.Y (nx16233), .A0 (camera_module_cache_ram_178__5), .A1 (
             nx35456), .S0 (nx34950)) ;
    dffr camera_module_cache_reg_ram_162__5 (.Q (camera_module_cache_ram_162__5)
         , .QB (\$dummy [1609]), .D (nx16243), .CLK (clk), .R (rst)) ;
    mux21_ni ix16244 (.Y (nx16243), .A0 (camera_module_cache_ram_162__5), .A1 (
             nx35456), .S0 (nx34954)) ;
    aoi22 ix31338 (.Y (nx31337), .A0 (camera_module_cache_ram_194__5), .A1 (
          nx36316), .B0 (camera_module_cache_ram_210__5), .B1 (nx36356)) ;
    dffr camera_module_cache_reg_ram_194__5 (.Q (camera_module_cache_ram_194__5)
         , .QB (\$dummy [1610]), .D (nx16223), .CLK (clk), .R (rst)) ;
    mux21_ni ix16224 (.Y (nx16223), .A0 (camera_module_cache_ram_194__5), .A1 (
             nx35456), .S0 (nx34946)) ;
    dffr camera_module_cache_reg_ram_210__5 (.Q (camera_module_cache_ram_210__5)
         , .QB (\$dummy [1611]), .D (nx16213), .CLK (clk), .R (rst)) ;
    mux21_ni ix16214 (.Y (nx16213), .A0 (camera_module_cache_ram_210__5), .A1 (
             nx35456), .S0 (nx34942)) ;
    aoi22 ix31346 (.Y (nx31345), .A0 (camera_module_cache_ram_226__5), .A1 (
          nx36396), .B0 (camera_module_cache_ram_242__5), .B1 (nx36436)) ;
    dffr camera_module_cache_reg_ram_226__5 (.Q (camera_module_cache_ram_226__5)
         , .QB (\$dummy [1612]), .D (nx16203), .CLK (clk), .R (rst)) ;
    mux21_ni ix16204 (.Y (nx16203), .A0 (camera_module_cache_ram_226__5), .A1 (
             nx35456), .S0 (nx34938)) ;
    dffr camera_module_cache_reg_ram_242__5 (.Q (camera_module_cache_ram_242__5)
         , .QB (\$dummy [1613]), .D (nx16193), .CLK (clk), .R (rst)) ;
    mux21_ni ix16194 (.Y (nx16193), .A0 (camera_module_cache_ram_242__5), .A1 (
             nx35456), .S0 (nx34934)) ;
    oai21 ix31354 (.Y (nx31353), .A0 (nx19316), .A1 (nx19238), .B0 (nx36460)) ;
    nand04 ix19317 (.Y (nx19316), .A0 (nx31356), .A1 (nx31364), .A2 (nx31372), .A3 (
           nx31380)) ;
    aoi22 ix31357 (.Y (nx31356), .A0 (camera_module_cache_ram_3__5), .A1 (
          nx35836), .B0 (camera_module_cache_ram_19__5), .B1 (nx35876)) ;
    dffr camera_module_cache_reg_ram_3__5 (.Q (camera_module_cache_ram_3__5), .QB (
         \$dummy [1614]), .D (nx16183), .CLK (clk), .R (rst)) ;
    mux21_ni ix16184 (.Y (nx16183), .A0 (camera_module_cache_ram_3__5), .A1 (
             nx35456), .S0 (nx34924)) ;
    dffr camera_module_cache_reg_ram_19__5 (.Q (camera_module_cache_ram_19__5), 
         .QB (\$dummy [1615]), .D (nx16173), .CLK (clk), .R (rst)) ;
    mux21_ni ix16174 (.Y (nx16173), .A0 (camera_module_cache_ram_19__5), .A1 (
             nx35458), .S0 (nx34920)) ;
    aoi22 ix31365 (.Y (nx31364), .A0 (camera_module_cache_ram_35__5), .A1 (
          nx35916), .B0 (camera_module_cache_ram_51__5), .B1 (nx35956)) ;
    dffr camera_module_cache_reg_ram_35__5 (.Q (camera_module_cache_ram_35__5), 
         .QB (\$dummy [1616]), .D (nx16163), .CLK (clk), .R (rst)) ;
    mux21_ni ix16164 (.Y (nx16163), .A0 (camera_module_cache_ram_35__5), .A1 (
             nx35458), .S0 (nx34916)) ;
    dffr camera_module_cache_reg_ram_51__5 (.Q (camera_module_cache_ram_51__5), 
         .QB (\$dummy [1617]), .D (nx16153), .CLK (clk), .R (rst)) ;
    mux21_ni ix16154 (.Y (nx16153), .A0 (camera_module_cache_ram_51__5), .A1 (
             nx35458), .S0 (nx34912)) ;
    aoi22 ix31373 (.Y (nx31372), .A0 (camera_module_cache_ram_67__5), .A1 (
          nx35996), .B0 (camera_module_cache_ram_83__5), .B1 (nx36036)) ;
    dffr camera_module_cache_reg_ram_67__5 (.Q (camera_module_cache_ram_67__5), 
         .QB (\$dummy [1618]), .D (nx16143), .CLK (clk), .R (rst)) ;
    mux21_ni ix16144 (.Y (nx16143), .A0 (camera_module_cache_ram_67__5), .A1 (
             nx35458), .S0 (nx34908)) ;
    dffr camera_module_cache_reg_ram_83__5 (.Q (camera_module_cache_ram_83__5), 
         .QB (\$dummy [1619]), .D (nx16133), .CLK (clk), .R (rst)) ;
    mux21_ni ix16134 (.Y (nx16133), .A0 (camera_module_cache_ram_83__5), .A1 (
             nx35458), .S0 (nx34904)) ;
    aoi22 ix31381 (.Y (nx31380), .A0 (camera_module_cache_ram_115__5), .A1 (
          nx36076), .B0 (camera_module_cache_ram_99__5), .B1 (nx36116)) ;
    dffr camera_module_cache_reg_ram_115__5 (.Q (camera_module_cache_ram_115__5)
         , .QB (\$dummy [1620]), .D (nx16113), .CLK (clk), .R (rst)) ;
    mux21_ni ix16114 (.Y (nx16113), .A0 (camera_module_cache_ram_115__5), .A1 (
             nx35458), .S0 (nx34896)) ;
    dffr camera_module_cache_reg_ram_99__5 (.Q (camera_module_cache_ram_99__5), 
         .QB (\$dummy [1621]), .D (nx16123), .CLK (clk), .R (rst)) ;
    mux21_ni ix16124 (.Y (nx16123), .A0 (camera_module_cache_ram_99__5), .A1 (
             nx35458), .S0 (nx34900)) ;
    nand04 ix19239 (.Y (nx19238), .A0 (nx31389), .A1 (nx31397), .A2 (nx31405), .A3 (
           nx31413)) ;
    aoi22 ix31390 (.Y (nx31389), .A0 (camera_module_cache_ram_131__5), .A1 (
          nx36156), .B0 (camera_module_cache_ram_147__5), .B1 (nx36196)) ;
    dffr camera_module_cache_reg_ram_131__5 (.Q (camera_module_cache_ram_131__5)
         , .QB (\$dummy [1622]), .D (nx16103), .CLK (clk), .R (rst)) ;
    mux21_ni ix16104 (.Y (nx16103), .A0 (camera_module_cache_ram_131__5), .A1 (
             nx35460), .S0 (nx34892)) ;
    dffr camera_module_cache_reg_ram_147__5 (.Q (camera_module_cache_ram_147__5)
         , .QB (\$dummy [1623]), .D (nx16093), .CLK (clk), .R (rst)) ;
    mux21_ni ix16094 (.Y (nx16093), .A0 (camera_module_cache_ram_147__5), .A1 (
             nx35460), .S0 (nx34888)) ;
    aoi22 ix31398 (.Y (nx31397), .A0 (camera_module_cache_ram_179__5), .A1 (
          nx36236), .B0 (camera_module_cache_ram_163__5), .B1 (nx36276)) ;
    dffr camera_module_cache_reg_ram_179__5 (.Q (camera_module_cache_ram_179__5)
         , .QB (\$dummy [1624]), .D (nx16073), .CLK (clk), .R (rst)) ;
    mux21_ni ix16074 (.Y (nx16073), .A0 (camera_module_cache_ram_179__5), .A1 (
             nx35460), .S0 (nx34880)) ;
    dffr camera_module_cache_reg_ram_163__5 (.Q (camera_module_cache_ram_163__5)
         , .QB (\$dummy [1625]), .D (nx16083), .CLK (clk), .R (rst)) ;
    mux21_ni ix16084 (.Y (nx16083), .A0 (camera_module_cache_ram_163__5), .A1 (
             nx35460), .S0 (nx34884)) ;
    aoi22 ix31406 (.Y (nx31405), .A0 (camera_module_cache_ram_195__5), .A1 (
          nx36316), .B0 (camera_module_cache_ram_211__5), .B1 (nx36356)) ;
    dffr camera_module_cache_reg_ram_195__5 (.Q (camera_module_cache_ram_195__5)
         , .QB (\$dummy [1626]), .D (nx16063), .CLK (clk), .R (rst)) ;
    mux21_ni ix16064 (.Y (nx16063), .A0 (camera_module_cache_ram_195__5), .A1 (
             nx35460), .S0 (nx34876)) ;
    dffr camera_module_cache_reg_ram_211__5 (.Q (camera_module_cache_ram_211__5)
         , .QB (\$dummy [1627]), .D (nx16053), .CLK (clk), .R (rst)) ;
    mux21_ni ix16054 (.Y (nx16053), .A0 (camera_module_cache_ram_211__5), .A1 (
             nx35460), .S0 (nx34872)) ;
    aoi22 ix31414 (.Y (nx31413), .A0 (camera_module_cache_ram_227__5), .A1 (
          nx36396), .B0 (camera_module_cache_ram_243__5), .B1 (nx36436)) ;
    dffr camera_module_cache_reg_ram_227__5 (.Q (camera_module_cache_ram_227__5)
         , .QB (\$dummy [1628]), .D (nx16043), .CLK (clk), .R (rst)) ;
    mux21_ni ix16044 (.Y (nx16043), .A0 (camera_module_cache_ram_227__5), .A1 (
             nx35460), .S0 (nx34868)) ;
    dffr camera_module_cache_reg_ram_243__5 (.Q (camera_module_cache_ram_243__5)
         , .QB (\$dummy [1629]), .D (nx16033), .CLK (clk), .R (rst)) ;
    mux21_ni ix16034 (.Y (nx16033), .A0 (camera_module_cache_ram_243__5), .A1 (
             nx35462), .S0 (nx34864)) ;
    nand04 ix19161 (.Y (nx19160), .A0 (nx31422), .A1 (nx31490), .A2 (nx31558), .A3 (
           nx31626)) ;
    oai21 ix31423 (.Y (nx31422), .A0 (nx19150), .A1 (nx19072), .B0 (nx36464)) ;
    nand04 ix19151 (.Y (nx19150), .A0 (nx31425), .A1 (nx31433), .A2 (nx31441), .A3 (
           nx31449)) ;
    aoi22 ix31426 (.Y (nx31425), .A0 (camera_module_cache_ram_4__5), .A1 (
          nx35836), .B0 (camera_module_cache_ram_20__5), .B1 (nx35876)) ;
    dffr camera_module_cache_reg_ram_4__5 (.Q (camera_module_cache_ram_4__5), .QB (
         \$dummy [1630]), .D (nx16023), .CLK (clk), .R (rst)) ;
    mux21_ni ix16024 (.Y (nx16023), .A0 (camera_module_cache_ram_4__5), .A1 (
             nx35462), .S0 (nx34854)) ;
    dffr camera_module_cache_reg_ram_20__5 (.Q (camera_module_cache_ram_20__5), 
         .QB (\$dummy [1631]), .D (nx16013), .CLK (clk), .R (rst)) ;
    mux21_ni ix16014 (.Y (nx16013), .A0 (camera_module_cache_ram_20__5), .A1 (
             nx35462), .S0 (nx34850)) ;
    aoi22 ix31434 (.Y (nx31433), .A0 (camera_module_cache_ram_36__5), .A1 (
          nx35916), .B0 (camera_module_cache_ram_52__5), .B1 (nx35956)) ;
    dffr camera_module_cache_reg_ram_36__5 (.Q (camera_module_cache_ram_36__5), 
         .QB (\$dummy [1632]), .D (nx16003), .CLK (clk), .R (rst)) ;
    mux21_ni ix16004 (.Y (nx16003), .A0 (camera_module_cache_ram_36__5), .A1 (
             nx35462), .S0 (nx34846)) ;
    dffr camera_module_cache_reg_ram_52__5 (.Q (camera_module_cache_ram_52__5), 
         .QB (\$dummy [1633]), .D (nx15993), .CLK (clk), .R (rst)) ;
    mux21_ni ix15994 (.Y (nx15993), .A0 (camera_module_cache_ram_52__5), .A1 (
             nx35462), .S0 (nx34842)) ;
    aoi22 ix31442 (.Y (nx31441), .A0 (camera_module_cache_ram_68__5), .A1 (
          nx35996), .B0 (camera_module_cache_ram_84__5), .B1 (nx36036)) ;
    dffr camera_module_cache_reg_ram_68__5 (.Q (camera_module_cache_ram_68__5), 
         .QB (\$dummy [1634]), .D (nx15983), .CLK (clk), .R (rst)) ;
    mux21_ni ix15984 (.Y (nx15983), .A0 (camera_module_cache_ram_68__5), .A1 (
             nx35462), .S0 (nx34838)) ;
    dffr camera_module_cache_reg_ram_84__5 (.Q (camera_module_cache_ram_84__5), 
         .QB (\$dummy [1635]), .D (nx15973), .CLK (clk), .R (rst)) ;
    mux21_ni ix15974 (.Y (nx15973), .A0 (camera_module_cache_ram_84__5), .A1 (
             nx35462), .S0 (nx34834)) ;
    aoi22 ix31450 (.Y (nx31449), .A0 (camera_module_cache_ram_116__5), .A1 (
          nx36076), .B0 (camera_module_cache_ram_100__5), .B1 (nx36116)) ;
    dffr camera_module_cache_reg_ram_116__5 (.Q (camera_module_cache_ram_116__5)
         , .QB (\$dummy [1636]), .D (nx15953), .CLK (clk), .R (rst)) ;
    mux21_ni ix15954 (.Y (nx15953), .A0 (camera_module_cache_ram_116__5), .A1 (
             nx35464), .S0 (nx34826)) ;
    dffr camera_module_cache_reg_ram_100__5 (.Q (camera_module_cache_ram_100__5)
         , .QB (\$dummy [1637]), .D (nx15963), .CLK (clk), .R (rst)) ;
    mux21_ni ix15964 (.Y (nx15963), .A0 (camera_module_cache_ram_100__5), .A1 (
             nx35464), .S0 (nx34830)) ;
    nand04 ix19073 (.Y (nx19072), .A0 (nx31458), .A1 (nx31466), .A2 (nx31474), .A3 (
           nx31482)) ;
    aoi22 ix31459 (.Y (nx31458), .A0 (camera_module_cache_ram_132__5), .A1 (
          nx36156), .B0 (camera_module_cache_ram_148__5), .B1 (nx36196)) ;
    dffr camera_module_cache_reg_ram_132__5 (.Q (camera_module_cache_ram_132__5)
         , .QB (\$dummy [1638]), .D (nx15943), .CLK (clk), .R (rst)) ;
    mux21_ni ix15944 (.Y (nx15943), .A0 (camera_module_cache_ram_132__5), .A1 (
             nx35464), .S0 (nx34822)) ;
    dffr camera_module_cache_reg_ram_148__5 (.Q (camera_module_cache_ram_148__5)
         , .QB (\$dummy [1639]), .D (nx15933), .CLK (clk), .R (rst)) ;
    mux21_ni ix15934 (.Y (nx15933), .A0 (camera_module_cache_ram_148__5), .A1 (
             nx35464), .S0 (nx34818)) ;
    aoi22 ix31467 (.Y (nx31466), .A0 (camera_module_cache_ram_180__5), .A1 (
          nx36236), .B0 (camera_module_cache_ram_164__5), .B1 (nx36276)) ;
    dffr camera_module_cache_reg_ram_180__5 (.Q (camera_module_cache_ram_180__5)
         , .QB (\$dummy [1640]), .D (nx15913), .CLK (clk), .R (rst)) ;
    mux21_ni ix15914 (.Y (nx15913), .A0 (camera_module_cache_ram_180__5), .A1 (
             nx35464), .S0 (nx34810)) ;
    dffr camera_module_cache_reg_ram_164__5 (.Q (camera_module_cache_ram_164__5)
         , .QB (\$dummy [1641]), .D (nx15923), .CLK (clk), .R (rst)) ;
    mux21_ni ix15924 (.Y (nx15923), .A0 (camera_module_cache_ram_164__5), .A1 (
             nx35464), .S0 (nx34814)) ;
    aoi22 ix31475 (.Y (nx31474), .A0 (camera_module_cache_ram_196__5), .A1 (
          nx36316), .B0 (camera_module_cache_ram_212__5), .B1 (nx36356)) ;
    dffr camera_module_cache_reg_ram_196__5 (.Q (camera_module_cache_ram_196__5)
         , .QB (\$dummy [1642]), .D (nx15903), .CLK (clk), .R (rst)) ;
    mux21_ni ix15904 (.Y (nx15903), .A0 (camera_module_cache_ram_196__5), .A1 (
             nx35464), .S0 (nx34806)) ;
    dffr camera_module_cache_reg_ram_212__5 (.Q (camera_module_cache_ram_212__5)
         , .QB (\$dummy [1643]), .D (nx15893), .CLK (clk), .R (rst)) ;
    mux21_ni ix15894 (.Y (nx15893), .A0 (camera_module_cache_ram_212__5), .A1 (
             nx35466), .S0 (nx34802)) ;
    aoi22 ix31483 (.Y (nx31482), .A0 (camera_module_cache_ram_228__5), .A1 (
          nx36396), .B0 (camera_module_cache_ram_244__5), .B1 (nx36436)) ;
    dffr camera_module_cache_reg_ram_228__5 (.Q (camera_module_cache_ram_228__5)
         , .QB (\$dummy [1644]), .D (nx15883), .CLK (clk), .R (rst)) ;
    mux21_ni ix15884 (.Y (nx15883), .A0 (camera_module_cache_ram_228__5), .A1 (
             nx35466), .S0 (nx34798)) ;
    dffr camera_module_cache_reg_ram_244__5 (.Q (camera_module_cache_ram_244__5)
         , .QB (\$dummy [1645]), .D (nx15873), .CLK (clk), .R (rst)) ;
    mux21_ni ix15874 (.Y (nx15873), .A0 (camera_module_cache_ram_244__5), .A1 (
             nx35466), .S0 (nx34794)) ;
    oai21 ix31491 (.Y (nx31490), .A0 (nx18988), .A1 (nx18910), .B0 (nx36468)) ;
    nand04 ix18989 (.Y (nx18988), .A0 (nx31493), .A1 (nx31501), .A2 (nx31509), .A3 (
           nx31517)) ;
    aoi22 ix31494 (.Y (nx31493), .A0 (camera_module_cache_ram_5__5), .A1 (
          nx35838), .B0 (camera_module_cache_ram_21__5), .B1 (nx35878)) ;
    dffr camera_module_cache_reg_ram_5__5 (.Q (camera_module_cache_ram_5__5), .QB (
         \$dummy [1646]), .D (nx15863), .CLK (clk), .R (rst)) ;
    mux21_ni ix15864 (.Y (nx15863), .A0 (camera_module_cache_ram_5__5), .A1 (
             nx35466), .S0 (nx34784)) ;
    dffr camera_module_cache_reg_ram_21__5 (.Q (camera_module_cache_ram_21__5), 
         .QB (\$dummy [1647]), .D (nx15853), .CLK (clk), .R (rst)) ;
    mux21_ni ix15854 (.Y (nx15853), .A0 (camera_module_cache_ram_21__5), .A1 (
             nx35466), .S0 (nx34780)) ;
    aoi22 ix31502 (.Y (nx31501), .A0 (camera_module_cache_ram_37__5), .A1 (
          nx35918), .B0 (camera_module_cache_ram_53__5), .B1 (nx35958)) ;
    dffr camera_module_cache_reg_ram_37__5 (.Q (camera_module_cache_ram_37__5), 
         .QB (\$dummy [1648]), .D (nx15843), .CLK (clk), .R (rst)) ;
    mux21_ni ix15844 (.Y (nx15843), .A0 (camera_module_cache_ram_37__5), .A1 (
             nx35466), .S0 (nx34776)) ;
    dffr camera_module_cache_reg_ram_53__5 (.Q (camera_module_cache_ram_53__5), 
         .QB (\$dummy [1649]), .D (nx15833), .CLK (clk), .R (rst)) ;
    mux21_ni ix15834 (.Y (nx15833), .A0 (camera_module_cache_ram_53__5), .A1 (
             nx35466), .S0 (nx34772)) ;
    aoi22 ix31510 (.Y (nx31509), .A0 (camera_module_cache_ram_69__5), .A1 (
          nx35998), .B0 (camera_module_cache_ram_85__5), .B1 (nx36038)) ;
    dffr camera_module_cache_reg_ram_69__5 (.Q (camera_module_cache_ram_69__5), 
         .QB (\$dummy [1650]), .D (nx15823), .CLK (clk), .R (rst)) ;
    mux21_ni ix15824 (.Y (nx15823), .A0 (camera_module_cache_ram_69__5), .A1 (
             nx35468), .S0 (nx34768)) ;
    dffr camera_module_cache_reg_ram_85__5 (.Q (camera_module_cache_ram_85__5), 
         .QB (\$dummy [1651]), .D (nx15813), .CLK (clk), .R (rst)) ;
    mux21_ni ix15814 (.Y (nx15813), .A0 (camera_module_cache_ram_85__5), .A1 (
             nx35468), .S0 (nx34764)) ;
    aoi22 ix31518 (.Y (nx31517), .A0 (camera_module_cache_ram_117__5), .A1 (
          nx36078), .B0 (camera_module_cache_ram_101__5), .B1 (nx36118)) ;
    dffr camera_module_cache_reg_ram_117__5 (.Q (camera_module_cache_ram_117__5)
         , .QB (\$dummy [1652]), .D (nx15793), .CLK (clk), .R (rst)) ;
    mux21_ni ix15794 (.Y (nx15793), .A0 (camera_module_cache_ram_117__5), .A1 (
             nx35468), .S0 (nx34756)) ;
    dffr camera_module_cache_reg_ram_101__5 (.Q (camera_module_cache_ram_101__5)
         , .QB (\$dummy [1653]), .D (nx15803), .CLK (clk), .R (rst)) ;
    mux21_ni ix15804 (.Y (nx15803), .A0 (camera_module_cache_ram_101__5), .A1 (
             nx35468), .S0 (nx34760)) ;
    nand04 ix18911 (.Y (nx18910), .A0 (nx31526), .A1 (nx31534), .A2 (nx31542), .A3 (
           nx31550)) ;
    aoi22 ix31527 (.Y (nx31526), .A0 (camera_module_cache_ram_133__5), .A1 (
          nx36158), .B0 (camera_module_cache_ram_149__5), .B1 (nx36198)) ;
    dffr camera_module_cache_reg_ram_133__5 (.Q (camera_module_cache_ram_133__5)
         , .QB (\$dummy [1654]), .D (nx15783), .CLK (clk), .R (rst)) ;
    mux21_ni ix15784 (.Y (nx15783), .A0 (camera_module_cache_ram_133__5), .A1 (
             nx35468), .S0 (nx34752)) ;
    dffr camera_module_cache_reg_ram_149__5 (.Q (camera_module_cache_ram_149__5)
         , .QB (\$dummy [1655]), .D (nx15773), .CLK (clk), .R (rst)) ;
    mux21_ni ix15774 (.Y (nx15773), .A0 (camera_module_cache_ram_149__5), .A1 (
             nx35468), .S0 (nx34748)) ;
    aoi22 ix31535 (.Y (nx31534), .A0 (camera_module_cache_ram_181__5), .A1 (
          nx36238), .B0 (camera_module_cache_ram_165__5), .B1 (nx36278)) ;
    dffr camera_module_cache_reg_ram_181__5 (.Q (camera_module_cache_ram_181__5)
         , .QB (\$dummy [1656]), .D (nx15753), .CLK (clk), .R (rst)) ;
    mux21_ni ix15754 (.Y (nx15753), .A0 (camera_module_cache_ram_181__5), .A1 (
             nx35468), .S0 (nx34740)) ;
    dffr camera_module_cache_reg_ram_165__5 (.Q (camera_module_cache_ram_165__5)
         , .QB (\$dummy [1657]), .D (nx15763), .CLK (clk), .R (rst)) ;
    mux21_ni ix15764 (.Y (nx15763), .A0 (camera_module_cache_ram_165__5), .A1 (
             nx35470), .S0 (nx34744)) ;
    aoi22 ix31543 (.Y (nx31542), .A0 (camera_module_cache_ram_197__5), .A1 (
          nx36318), .B0 (camera_module_cache_ram_213__5), .B1 (nx36358)) ;
    dffr camera_module_cache_reg_ram_197__5 (.Q (camera_module_cache_ram_197__5)
         , .QB (\$dummy [1658]), .D (nx15743), .CLK (clk), .R (rst)) ;
    mux21_ni ix15744 (.Y (nx15743), .A0 (camera_module_cache_ram_197__5), .A1 (
             nx35470), .S0 (nx34736)) ;
    dffr camera_module_cache_reg_ram_213__5 (.Q (camera_module_cache_ram_213__5)
         , .QB (\$dummy [1659]), .D (nx15733), .CLK (clk), .R (rst)) ;
    mux21_ni ix15734 (.Y (nx15733), .A0 (camera_module_cache_ram_213__5), .A1 (
             nx35470), .S0 (nx34732)) ;
    aoi22 ix31551 (.Y (nx31550), .A0 (camera_module_cache_ram_229__5), .A1 (
          nx36398), .B0 (camera_module_cache_ram_245__5), .B1 (nx36438)) ;
    dffr camera_module_cache_reg_ram_229__5 (.Q (camera_module_cache_ram_229__5)
         , .QB (\$dummy [1660]), .D (nx15723), .CLK (clk), .R (rst)) ;
    mux21_ni ix15724 (.Y (nx15723), .A0 (camera_module_cache_ram_229__5), .A1 (
             nx35470), .S0 (nx34728)) ;
    dffr camera_module_cache_reg_ram_245__5 (.Q (camera_module_cache_ram_245__5)
         , .QB (\$dummy [1661]), .D (nx15713), .CLK (clk), .R (rst)) ;
    mux21_ni ix15714 (.Y (nx15713), .A0 (camera_module_cache_ram_245__5), .A1 (
             nx35470), .S0 (nx34724)) ;
    oai21 ix31559 (.Y (nx31558), .A0 (nx18824), .A1 (nx18746), .B0 (nx36472)) ;
    nand04 ix18825 (.Y (nx18824), .A0 (nx31561), .A1 (nx31569), .A2 (nx31577), .A3 (
           nx31585)) ;
    aoi22 ix31562 (.Y (nx31561), .A0 (camera_module_cache_ram_6__5), .A1 (
          nx35838), .B0 (camera_module_cache_ram_22__5), .B1 (nx35878)) ;
    dffr camera_module_cache_reg_ram_6__5 (.Q (camera_module_cache_ram_6__5), .QB (
         \$dummy [1662]), .D (nx15703), .CLK (clk), .R (rst)) ;
    mux21_ni ix15704 (.Y (nx15703), .A0 (camera_module_cache_ram_6__5), .A1 (
             nx35470), .S0 (nx34714)) ;
    dffr camera_module_cache_reg_ram_22__5 (.Q (camera_module_cache_ram_22__5), 
         .QB (\$dummy [1663]), .D (nx15693), .CLK (clk), .R (rst)) ;
    mux21_ni ix15694 (.Y (nx15693), .A0 (camera_module_cache_ram_22__5), .A1 (
             nx35470), .S0 (nx34710)) ;
    aoi22 ix31570 (.Y (nx31569), .A0 (camera_module_cache_ram_38__5), .A1 (
          nx35918), .B0 (camera_module_cache_ram_54__5), .B1 (nx35958)) ;
    dffr camera_module_cache_reg_ram_38__5 (.Q (camera_module_cache_ram_38__5), 
         .QB (\$dummy [1664]), .D (nx15683), .CLK (clk), .R (rst)) ;
    mux21_ni ix15684 (.Y (nx15683), .A0 (camera_module_cache_ram_38__5), .A1 (
             nx35472), .S0 (nx34706)) ;
    dffr camera_module_cache_reg_ram_54__5 (.Q (camera_module_cache_ram_54__5), 
         .QB (\$dummy [1665]), .D (nx15673), .CLK (clk), .R (rst)) ;
    mux21_ni ix15674 (.Y (nx15673), .A0 (camera_module_cache_ram_54__5), .A1 (
             nx35472), .S0 (nx34702)) ;
    aoi22 ix31578 (.Y (nx31577), .A0 (camera_module_cache_ram_70__5), .A1 (
          nx35998), .B0 (camera_module_cache_ram_86__5), .B1 (nx36038)) ;
    dffr camera_module_cache_reg_ram_70__5 (.Q (camera_module_cache_ram_70__5), 
         .QB (\$dummy [1666]), .D (nx15663), .CLK (clk), .R (rst)) ;
    mux21_ni ix15664 (.Y (nx15663), .A0 (camera_module_cache_ram_70__5), .A1 (
             nx35472), .S0 (nx34698)) ;
    dffr camera_module_cache_reg_ram_86__5 (.Q (camera_module_cache_ram_86__5), 
         .QB (\$dummy [1667]), .D (nx15653), .CLK (clk), .R (rst)) ;
    mux21_ni ix15654 (.Y (nx15653), .A0 (camera_module_cache_ram_86__5), .A1 (
             nx35472), .S0 (nx34694)) ;
    aoi22 ix31586 (.Y (nx31585), .A0 (camera_module_cache_ram_118__5), .A1 (
          nx36078), .B0 (camera_module_cache_ram_102__5), .B1 (nx36118)) ;
    dffr camera_module_cache_reg_ram_118__5 (.Q (camera_module_cache_ram_118__5)
         , .QB (\$dummy [1668]), .D (nx15633), .CLK (clk), .R (rst)) ;
    mux21_ni ix15634 (.Y (nx15633), .A0 (camera_module_cache_ram_118__5), .A1 (
             nx35472), .S0 (nx34686)) ;
    dffr camera_module_cache_reg_ram_102__5 (.Q (camera_module_cache_ram_102__5)
         , .QB (\$dummy [1669]), .D (nx15643), .CLK (clk), .R (rst)) ;
    mux21_ni ix15644 (.Y (nx15643), .A0 (camera_module_cache_ram_102__5), .A1 (
             nx35472), .S0 (nx34690)) ;
    nand04 ix18747 (.Y (nx18746), .A0 (nx31594), .A1 (nx31602), .A2 (nx31610), .A3 (
           nx31618)) ;
    aoi22 ix31595 (.Y (nx31594), .A0 (camera_module_cache_ram_134__5), .A1 (
          nx36158), .B0 (camera_module_cache_ram_150__5), .B1 (nx36198)) ;
    dffr camera_module_cache_reg_ram_134__5 (.Q (camera_module_cache_ram_134__5)
         , .QB (\$dummy [1670]), .D (nx15623), .CLK (clk), .R (rst)) ;
    mux21_ni ix15624 (.Y (nx15623), .A0 (camera_module_cache_ram_134__5), .A1 (
             nx35472), .S0 (nx34682)) ;
    dffr camera_module_cache_reg_ram_150__5 (.Q (camera_module_cache_ram_150__5)
         , .QB (\$dummy [1671]), .D (nx15613), .CLK (clk), .R (rst)) ;
    mux21_ni ix15614 (.Y (nx15613), .A0 (camera_module_cache_ram_150__5), .A1 (
             nx35474), .S0 (nx34678)) ;
    aoi22 ix31603 (.Y (nx31602), .A0 (camera_module_cache_ram_182__5), .A1 (
          nx36238), .B0 (camera_module_cache_ram_166__5), .B1 (nx36278)) ;
    dffr camera_module_cache_reg_ram_182__5 (.Q (camera_module_cache_ram_182__5)
         , .QB (\$dummy [1672]), .D (nx15593), .CLK (clk), .R (rst)) ;
    mux21_ni ix15594 (.Y (nx15593), .A0 (camera_module_cache_ram_182__5), .A1 (
             nx35474), .S0 (nx34670)) ;
    dffr camera_module_cache_reg_ram_166__5 (.Q (camera_module_cache_ram_166__5)
         , .QB (\$dummy [1673]), .D (nx15603), .CLK (clk), .R (rst)) ;
    mux21_ni ix15604 (.Y (nx15603), .A0 (camera_module_cache_ram_166__5), .A1 (
             nx35474), .S0 (nx34674)) ;
    aoi22 ix31611 (.Y (nx31610), .A0 (camera_module_cache_ram_198__5), .A1 (
          nx36318), .B0 (camera_module_cache_ram_214__5), .B1 (nx36358)) ;
    dffr camera_module_cache_reg_ram_198__5 (.Q (camera_module_cache_ram_198__5)
         , .QB (\$dummy [1674]), .D (nx15583), .CLK (clk), .R (rst)) ;
    mux21_ni ix15584 (.Y (nx15583), .A0 (camera_module_cache_ram_198__5), .A1 (
             nx35474), .S0 (nx34666)) ;
    dffr camera_module_cache_reg_ram_214__5 (.Q (camera_module_cache_ram_214__5)
         , .QB (\$dummy [1675]), .D (nx15573), .CLK (clk), .R (rst)) ;
    mux21_ni ix15574 (.Y (nx15573), .A0 (camera_module_cache_ram_214__5), .A1 (
             nx35474), .S0 (nx34662)) ;
    aoi22 ix31619 (.Y (nx31618), .A0 (camera_module_cache_ram_230__5), .A1 (
          nx36398), .B0 (camera_module_cache_ram_246__5), .B1 (nx36438)) ;
    dffr camera_module_cache_reg_ram_230__5 (.Q (camera_module_cache_ram_230__5)
         , .QB (\$dummy [1676]), .D (nx15563), .CLK (clk), .R (rst)) ;
    mux21_ni ix15564 (.Y (nx15563), .A0 (camera_module_cache_ram_230__5), .A1 (
             nx35474), .S0 (nx34658)) ;
    dffr camera_module_cache_reg_ram_246__5 (.Q (camera_module_cache_ram_246__5)
         , .QB (\$dummy [1677]), .D (nx15553), .CLK (clk), .R (rst)) ;
    mux21_ni ix15554 (.Y (nx15553), .A0 (camera_module_cache_ram_246__5), .A1 (
             nx35474), .S0 (nx34654)) ;
    oai21 ix31627 (.Y (nx31626), .A0 (nx18662), .A1 (nx18584), .B0 (nx36476)) ;
    nand04 ix18663 (.Y (nx18662), .A0 (nx31629), .A1 (nx31637), .A2 (nx31645), .A3 (
           nx31653)) ;
    aoi22 ix31630 (.Y (nx31629), .A0 (camera_module_cache_ram_7__5), .A1 (
          nx35838), .B0 (camera_module_cache_ram_23__5), .B1 (nx35878)) ;
    dffr camera_module_cache_reg_ram_7__5 (.Q (camera_module_cache_ram_7__5), .QB (
         \$dummy [1678]), .D (nx15543), .CLK (clk), .R (rst)) ;
    mux21_ni ix15544 (.Y (nx15543), .A0 (camera_module_cache_ram_7__5), .A1 (
             nx35476), .S0 (nx34644)) ;
    dffr camera_module_cache_reg_ram_23__5 (.Q (camera_module_cache_ram_23__5), 
         .QB (\$dummy [1679]), .D (nx15533), .CLK (clk), .R (rst)) ;
    mux21_ni ix15534 (.Y (nx15533), .A0 (camera_module_cache_ram_23__5), .A1 (
             nx35476), .S0 (nx34640)) ;
    aoi22 ix31638 (.Y (nx31637), .A0 (camera_module_cache_ram_39__5), .A1 (
          nx35918), .B0 (camera_module_cache_ram_55__5), .B1 (nx35958)) ;
    dffr camera_module_cache_reg_ram_39__5 (.Q (camera_module_cache_ram_39__5), 
         .QB (\$dummy [1680]), .D (nx15523), .CLK (clk), .R (rst)) ;
    mux21_ni ix15524 (.Y (nx15523), .A0 (camera_module_cache_ram_39__5), .A1 (
             nx35476), .S0 (nx34636)) ;
    dffr camera_module_cache_reg_ram_55__5 (.Q (camera_module_cache_ram_55__5), 
         .QB (\$dummy [1681]), .D (nx15513), .CLK (clk), .R (rst)) ;
    mux21_ni ix15514 (.Y (nx15513), .A0 (camera_module_cache_ram_55__5), .A1 (
             nx35476), .S0 (nx34632)) ;
    aoi22 ix31646 (.Y (nx31645), .A0 (camera_module_cache_ram_71__5), .A1 (
          nx35998), .B0 (camera_module_cache_ram_87__5), .B1 (nx36038)) ;
    dffr camera_module_cache_reg_ram_71__5 (.Q (camera_module_cache_ram_71__5), 
         .QB (\$dummy [1682]), .D (nx15503), .CLK (clk), .R (rst)) ;
    mux21_ni ix15504 (.Y (nx15503), .A0 (camera_module_cache_ram_71__5), .A1 (
             nx35476), .S0 (nx34628)) ;
    dffr camera_module_cache_reg_ram_87__5 (.Q (camera_module_cache_ram_87__5), 
         .QB (\$dummy [1683]), .D (nx15493), .CLK (clk), .R (rst)) ;
    mux21_ni ix15494 (.Y (nx15493), .A0 (camera_module_cache_ram_87__5), .A1 (
             nx35476), .S0 (nx34624)) ;
    aoi22 ix31654 (.Y (nx31653), .A0 (camera_module_cache_ram_119__5), .A1 (
          nx36078), .B0 (camera_module_cache_ram_103__5), .B1 (nx36118)) ;
    dffr camera_module_cache_reg_ram_119__5 (.Q (camera_module_cache_ram_119__5)
         , .QB (\$dummy [1684]), .D (nx15473), .CLK (clk), .R (rst)) ;
    mux21_ni ix15474 (.Y (nx15473), .A0 (camera_module_cache_ram_119__5), .A1 (
             nx35476), .S0 (nx34616)) ;
    dffr camera_module_cache_reg_ram_103__5 (.Q (camera_module_cache_ram_103__5)
         , .QB (\$dummy [1685]), .D (nx15483), .CLK (clk), .R (rst)) ;
    mux21_ni ix15484 (.Y (nx15483), .A0 (camera_module_cache_ram_103__5), .A1 (
             nx35478), .S0 (nx34620)) ;
    nand04 ix18585 (.Y (nx18584), .A0 (nx31662), .A1 (nx31670), .A2 (nx31678), .A3 (
           nx31686)) ;
    aoi22 ix31663 (.Y (nx31662), .A0 (camera_module_cache_ram_135__5), .A1 (
          nx36158), .B0 (camera_module_cache_ram_151__5), .B1 (nx36198)) ;
    dffr camera_module_cache_reg_ram_135__5 (.Q (camera_module_cache_ram_135__5)
         , .QB (\$dummy [1686]), .D (nx15463), .CLK (clk), .R (rst)) ;
    mux21_ni ix15464 (.Y (nx15463), .A0 (camera_module_cache_ram_135__5), .A1 (
             nx35478), .S0 (nx34612)) ;
    dffr camera_module_cache_reg_ram_151__5 (.Q (camera_module_cache_ram_151__5)
         , .QB (\$dummy [1687]), .D (nx15453), .CLK (clk), .R (rst)) ;
    mux21_ni ix15454 (.Y (nx15453), .A0 (camera_module_cache_ram_151__5), .A1 (
             nx35478), .S0 (nx34608)) ;
    aoi22 ix31671 (.Y (nx31670), .A0 (camera_module_cache_ram_183__5), .A1 (
          nx36238), .B0 (camera_module_cache_ram_167__5), .B1 (nx36278)) ;
    dffr camera_module_cache_reg_ram_183__5 (.Q (camera_module_cache_ram_183__5)
         , .QB (\$dummy [1688]), .D (nx15433), .CLK (clk), .R (rst)) ;
    mux21_ni ix15434 (.Y (nx15433), .A0 (camera_module_cache_ram_183__5), .A1 (
             nx35478), .S0 (nx34600)) ;
    dffr camera_module_cache_reg_ram_167__5 (.Q (camera_module_cache_ram_167__5)
         , .QB (\$dummy [1689]), .D (nx15443), .CLK (clk), .R (rst)) ;
    mux21_ni ix15444 (.Y (nx15443), .A0 (camera_module_cache_ram_167__5), .A1 (
             nx35478), .S0 (nx34604)) ;
    aoi22 ix31679 (.Y (nx31678), .A0 (camera_module_cache_ram_199__5), .A1 (
          nx36318), .B0 (camera_module_cache_ram_215__5), .B1 (nx36358)) ;
    dffr camera_module_cache_reg_ram_199__5 (.Q (camera_module_cache_ram_199__5)
         , .QB (\$dummy [1690]), .D (nx15423), .CLK (clk), .R (rst)) ;
    mux21_ni ix15424 (.Y (nx15423), .A0 (camera_module_cache_ram_199__5), .A1 (
             nx35478), .S0 (nx34596)) ;
    dffr camera_module_cache_reg_ram_215__5 (.Q (camera_module_cache_ram_215__5)
         , .QB (\$dummy [1691]), .D (nx15413), .CLK (clk), .R (rst)) ;
    mux21_ni ix15414 (.Y (nx15413), .A0 (camera_module_cache_ram_215__5), .A1 (
             nx35478), .S0 (nx34592)) ;
    aoi22 ix31687 (.Y (nx31686), .A0 (camera_module_cache_ram_231__5), .A1 (
          nx36398), .B0 (camera_module_cache_ram_247__5), .B1 (nx36438)) ;
    dffr camera_module_cache_reg_ram_231__5 (.Q (camera_module_cache_ram_231__5)
         , .QB (\$dummy [1692]), .D (nx15403), .CLK (clk), .R (rst)) ;
    mux21_ni ix15404 (.Y (nx15403), .A0 (camera_module_cache_ram_231__5), .A1 (
             nx35480), .S0 (nx34588)) ;
    dffr camera_module_cache_reg_ram_247__5 (.Q (camera_module_cache_ram_247__5)
         , .QB (\$dummy [1693]), .D (nx15393), .CLK (clk), .R (rst)) ;
    mux21_ni ix15394 (.Y (nx15393), .A0 (camera_module_cache_ram_247__5), .A1 (
             nx35480), .S0 (nx34584)) ;
    nand04 ix18505 (.Y (nx18504), .A0 (nx31695), .A1 (nx31763), .A2 (nx31831), .A3 (
           nx31899)) ;
    oai21 ix31696 (.Y (nx31695), .A0 (nx18494), .A1 (nx18416), .B0 (nx36480)) ;
    nand04 ix18495 (.Y (nx18494), .A0 (nx31698), .A1 (nx31706), .A2 (nx31714), .A3 (
           nx31722)) ;
    aoi22 ix31699 (.Y (nx31698), .A0 (camera_module_cache_ram_8__5), .A1 (
          nx35838), .B0 (camera_module_cache_ram_24__5), .B1 (nx35878)) ;
    dffr camera_module_cache_reg_ram_8__5 (.Q (camera_module_cache_ram_8__5), .QB (
         \$dummy [1694]), .D (nx15383), .CLK (clk), .R (rst)) ;
    mux21_ni ix15384 (.Y (nx15383), .A0 (camera_module_cache_ram_8__5), .A1 (
             nx35480), .S0 (nx34574)) ;
    dffr camera_module_cache_reg_ram_24__5 (.Q (camera_module_cache_ram_24__5), 
         .QB (\$dummy [1695]), .D (nx15373), .CLK (clk), .R (rst)) ;
    mux21_ni ix15374 (.Y (nx15373), .A0 (camera_module_cache_ram_24__5), .A1 (
             nx35480), .S0 (nx34570)) ;
    aoi22 ix31707 (.Y (nx31706), .A0 (camera_module_cache_ram_40__5), .A1 (
          nx35918), .B0 (camera_module_cache_ram_56__5), .B1 (nx35958)) ;
    dffr camera_module_cache_reg_ram_40__5 (.Q (camera_module_cache_ram_40__5), 
         .QB (\$dummy [1696]), .D (nx15363), .CLK (clk), .R (rst)) ;
    mux21_ni ix15364 (.Y (nx15363), .A0 (camera_module_cache_ram_40__5), .A1 (
             nx35480), .S0 (nx34566)) ;
    dffr camera_module_cache_reg_ram_56__5 (.Q (camera_module_cache_ram_56__5), 
         .QB (\$dummy [1697]), .D (nx15353), .CLK (clk), .R (rst)) ;
    mux21_ni ix15354 (.Y (nx15353), .A0 (camera_module_cache_ram_56__5), .A1 (
             nx35480), .S0 (nx34562)) ;
    aoi22 ix31715 (.Y (nx31714), .A0 (camera_module_cache_ram_72__5), .A1 (
          nx35998), .B0 (camera_module_cache_ram_88__5), .B1 (nx36038)) ;
    dffr camera_module_cache_reg_ram_72__5 (.Q (camera_module_cache_ram_72__5), 
         .QB (\$dummy [1698]), .D (nx15343), .CLK (clk), .R (rst)) ;
    mux21_ni ix15344 (.Y (nx15343), .A0 (camera_module_cache_ram_72__5), .A1 (
             nx35480), .S0 (nx34558)) ;
    dffr camera_module_cache_reg_ram_88__5 (.Q (camera_module_cache_ram_88__5), 
         .QB (\$dummy [1699]), .D (nx15333), .CLK (clk), .R (rst)) ;
    mux21_ni ix15334 (.Y (nx15333), .A0 (camera_module_cache_ram_88__5), .A1 (
             nx35482), .S0 (nx34554)) ;
    aoi22 ix31723 (.Y (nx31722), .A0 (camera_module_cache_ram_120__5), .A1 (
          nx36078), .B0 (camera_module_cache_ram_104__5), .B1 (nx36118)) ;
    dffr camera_module_cache_reg_ram_120__5 (.Q (camera_module_cache_ram_120__5)
         , .QB (\$dummy [1700]), .D (nx15313), .CLK (clk), .R (rst)) ;
    mux21_ni ix15314 (.Y (nx15313), .A0 (camera_module_cache_ram_120__5), .A1 (
             nx35482), .S0 (nx34546)) ;
    dffr camera_module_cache_reg_ram_104__5 (.Q (camera_module_cache_ram_104__5)
         , .QB (\$dummy [1701]), .D (nx15323), .CLK (clk), .R (rst)) ;
    mux21_ni ix15324 (.Y (nx15323), .A0 (camera_module_cache_ram_104__5), .A1 (
             nx35482), .S0 (nx34550)) ;
    nand04 ix18417 (.Y (nx18416), .A0 (nx31731), .A1 (nx31739), .A2 (nx31747), .A3 (
           nx31755)) ;
    aoi22 ix31732 (.Y (nx31731), .A0 (camera_module_cache_ram_136__5), .A1 (
          nx36158), .B0 (camera_module_cache_ram_152__5), .B1 (nx36198)) ;
    dffr camera_module_cache_reg_ram_136__5 (.Q (camera_module_cache_ram_136__5)
         , .QB (\$dummy [1702]), .D (nx15303), .CLK (clk), .R (rst)) ;
    mux21_ni ix15304 (.Y (nx15303), .A0 (camera_module_cache_ram_136__5), .A1 (
             nx35482), .S0 (nx34542)) ;
    dffr camera_module_cache_reg_ram_152__5 (.Q (camera_module_cache_ram_152__5)
         , .QB (\$dummy [1703]), .D (nx15293), .CLK (clk), .R (rst)) ;
    mux21_ni ix15294 (.Y (nx15293), .A0 (camera_module_cache_ram_152__5), .A1 (
             nx35482), .S0 (nx34538)) ;
    aoi22 ix31740 (.Y (nx31739), .A0 (camera_module_cache_ram_184__5), .A1 (
          nx36238), .B0 (camera_module_cache_ram_168__5), .B1 (nx36278)) ;
    dffr camera_module_cache_reg_ram_184__5 (.Q (camera_module_cache_ram_184__5)
         , .QB (\$dummy [1704]), .D (nx15273), .CLK (clk), .R (rst)) ;
    mux21_ni ix15274 (.Y (nx15273), .A0 (camera_module_cache_ram_184__5), .A1 (
             nx35482), .S0 (nx34530)) ;
    dffr camera_module_cache_reg_ram_168__5 (.Q (camera_module_cache_ram_168__5)
         , .QB (\$dummy [1705]), .D (nx15283), .CLK (clk), .R (rst)) ;
    mux21_ni ix15284 (.Y (nx15283), .A0 (camera_module_cache_ram_168__5), .A1 (
             nx35482), .S0 (nx34534)) ;
    aoi22 ix31748 (.Y (nx31747), .A0 (camera_module_cache_ram_200__5), .A1 (
          nx36318), .B0 (camera_module_cache_ram_216__5), .B1 (nx36358)) ;
    dffr camera_module_cache_reg_ram_200__5 (.Q (camera_module_cache_ram_200__5)
         , .QB (\$dummy [1706]), .D (nx15263), .CLK (clk), .R (rst)) ;
    mux21_ni ix15264 (.Y (nx15263), .A0 (camera_module_cache_ram_200__5), .A1 (
             nx35484), .S0 (nx34526)) ;
    dffr camera_module_cache_reg_ram_216__5 (.Q (camera_module_cache_ram_216__5)
         , .QB (\$dummy [1707]), .D (nx15253), .CLK (clk), .R (rst)) ;
    mux21_ni ix15254 (.Y (nx15253), .A0 (camera_module_cache_ram_216__5), .A1 (
             nx35484), .S0 (nx34522)) ;
    aoi22 ix31756 (.Y (nx31755), .A0 (camera_module_cache_ram_232__5), .A1 (
          nx36398), .B0 (camera_module_cache_ram_248__5), .B1 (nx36438)) ;
    dffr camera_module_cache_reg_ram_232__5 (.Q (camera_module_cache_ram_232__5)
         , .QB (\$dummy [1708]), .D (nx15243), .CLK (clk), .R (rst)) ;
    mux21_ni ix15244 (.Y (nx15243), .A0 (camera_module_cache_ram_232__5), .A1 (
             nx35484), .S0 (nx34518)) ;
    dffr camera_module_cache_reg_ram_248__5 (.Q (camera_module_cache_ram_248__5)
         , .QB (\$dummy [1709]), .D (nx15233), .CLK (clk), .R (rst)) ;
    mux21_ni ix15234 (.Y (nx15233), .A0 (camera_module_cache_ram_248__5), .A1 (
             nx35484), .S0 (nx34514)) ;
    oai21 ix31764 (.Y (nx31763), .A0 (nx18332), .A1 (nx18254), .B0 (nx36484)) ;
    nand04 ix18333 (.Y (nx18332), .A0 (nx31766), .A1 (nx31774), .A2 (nx31782), .A3 (
           nx31790)) ;
    aoi22 ix31767 (.Y (nx31766), .A0 (camera_module_cache_ram_9__5), .A1 (
          nx35838), .B0 (camera_module_cache_ram_25__5), .B1 (nx35878)) ;
    dffr camera_module_cache_reg_ram_9__5 (.Q (camera_module_cache_ram_9__5), .QB (
         \$dummy [1710]), .D (nx15223), .CLK (clk), .R (rst)) ;
    mux21_ni ix15224 (.Y (nx15223), .A0 (camera_module_cache_ram_9__5), .A1 (
             nx35484), .S0 (nx34504)) ;
    dffr camera_module_cache_reg_ram_25__5 (.Q (camera_module_cache_ram_25__5), 
         .QB (\$dummy [1711]), .D (nx15213), .CLK (clk), .R (rst)) ;
    mux21_ni ix15214 (.Y (nx15213), .A0 (camera_module_cache_ram_25__5), .A1 (
             nx35484), .S0 (nx34500)) ;
    aoi22 ix31775 (.Y (nx31774), .A0 (camera_module_cache_ram_41__5), .A1 (
          nx35918), .B0 (camera_module_cache_ram_57__5), .B1 (nx35958)) ;
    dffr camera_module_cache_reg_ram_41__5 (.Q (camera_module_cache_ram_41__5), 
         .QB (\$dummy [1712]), .D (nx15203), .CLK (clk), .R (rst)) ;
    mux21_ni ix15204 (.Y (nx15203), .A0 (camera_module_cache_ram_41__5), .A1 (
             nx35484), .S0 (nx34496)) ;
    dffr camera_module_cache_reg_ram_57__5 (.Q (camera_module_cache_ram_57__5), 
         .QB (\$dummy [1713]), .D (nx15193), .CLK (clk), .R (rst)) ;
    mux21_ni ix15194 (.Y (nx15193), .A0 (camera_module_cache_ram_57__5), .A1 (
             nx35486), .S0 (nx34492)) ;
    aoi22 ix31783 (.Y (nx31782), .A0 (camera_module_cache_ram_73__5), .A1 (
          nx35998), .B0 (camera_module_cache_ram_89__5), .B1 (nx36038)) ;
    dffr camera_module_cache_reg_ram_73__5 (.Q (camera_module_cache_ram_73__5), 
         .QB (\$dummy [1714]), .D (nx15183), .CLK (clk), .R (rst)) ;
    mux21_ni ix15184 (.Y (nx15183), .A0 (camera_module_cache_ram_73__5), .A1 (
             nx35486), .S0 (nx34488)) ;
    dffr camera_module_cache_reg_ram_89__5 (.Q (camera_module_cache_ram_89__5), 
         .QB (\$dummy [1715]), .D (nx15173), .CLK (clk), .R (rst)) ;
    mux21_ni ix15174 (.Y (nx15173), .A0 (camera_module_cache_ram_89__5), .A1 (
             nx35486), .S0 (nx34484)) ;
    aoi22 ix31791 (.Y (nx31790), .A0 (camera_module_cache_ram_121__5), .A1 (
          nx36078), .B0 (camera_module_cache_ram_105__5), .B1 (nx36118)) ;
    dffr camera_module_cache_reg_ram_121__5 (.Q (camera_module_cache_ram_121__5)
         , .QB (\$dummy [1716]), .D (nx15153), .CLK (clk), .R (rst)) ;
    mux21_ni ix15154 (.Y (nx15153), .A0 (camera_module_cache_ram_121__5), .A1 (
             nx35486), .S0 (nx34476)) ;
    dffr camera_module_cache_reg_ram_105__5 (.Q (camera_module_cache_ram_105__5)
         , .QB (\$dummy [1717]), .D (nx15163), .CLK (clk), .R (rst)) ;
    mux21_ni ix15164 (.Y (nx15163), .A0 (camera_module_cache_ram_105__5), .A1 (
             nx35486), .S0 (nx34480)) ;
    nand04 ix18255 (.Y (nx18254), .A0 (nx31799), .A1 (nx31807), .A2 (nx31815), .A3 (
           nx31823)) ;
    aoi22 ix31800 (.Y (nx31799), .A0 (camera_module_cache_ram_137__5), .A1 (
          nx36158), .B0 (camera_module_cache_ram_153__5), .B1 (nx36198)) ;
    dffr camera_module_cache_reg_ram_137__5 (.Q (camera_module_cache_ram_137__5)
         , .QB (\$dummy [1718]), .D (nx15143), .CLK (clk), .R (rst)) ;
    mux21_ni ix15144 (.Y (nx15143), .A0 (camera_module_cache_ram_137__5), .A1 (
             nx35486), .S0 (nx34472)) ;
    dffr camera_module_cache_reg_ram_153__5 (.Q (camera_module_cache_ram_153__5)
         , .QB (\$dummy [1719]), .D (nx15133), .CLK (clk), .R (rst)) ;
    mux21_ni ix15134 (.Y (nx15133), .A0 (camera_module_cache_ram_153__5), .A1 (
             nx35486), .S0 (nx34468)) ;
    aoi22 ix31808 (.Y (nx31807), .A0 (camera_module_cache_ram_185__5), .A1 (
          nx36238), .B0 (camera_module_cache_ram_169__5), .B1 (nx36278)) ;
    dffr camera_module_cache_reg_ram_185__5 (.Q (camera_module_cache_ram_185__5)
         , .QB (\$dummy [1720]), .D (nx15113), .CLK (clk), .R (rst)) ;
    mux21_ni ix15114 (.Y (nx15113), .A0 (camera_module_cache_ram_185__5), .A1 (
             nx35488), .S0 (nx34460)) ;
    dffr camera_module_cache_reg_ram_169__5 (.Q (camera_module_cache_ram_169__5)
         , .QB (\$dummy [1721]), .D (nx15123), .CLK (clk), .R (rst)) ;
    mux21_ni ix15124 (.Y (nx15123), .A0 (camera_module_cache_ram_169__5), .A1 (
             nx35488), .S0 (nx34464)) ;
    aoi22 ix31816 (.Y (nx31815), .A0 (camera_module_cache_ram_201__5), .A1 (
          nx36318), .B0 (camera_module_cache_ram_217__5), .B1 (nx36358)) ;
    dffr camera_module_cache_reg_ram_201__5 (.Q (camera_module_cache_ram_201__5)
         , .QB (\$dummy [1722]), .D (nx15103), .CLK (clk), .R (rst)) ;
    mux21_ni ix15104 (.Y (nx15103), .A0 (camera_module_cache_ram_201__5), .A1 (
             nx35488), .S0 (nx34456)) ;
    dffr camera_module_cache_reg_ram_217__5 (.Q (camera_module_cache_ram_217__5)
         , .QB (\$dummy [1723]), .D (nx15093), .CLK (clk), .R (rst)) ;
    mux21_ni ix15094 (.Y (nx15093), .A0 (camera_module_cache_ram_217__5), .A1 (
             nx35488), .S0 (nx34452)) ;
    aoi22 ix31824 (.Y (nx31823), .A0 (camera_module_cache_ram_233__5), .A1 (
          nx36398), .B0 (camera_module_cache_ram_249__5), .B1 (nx36438)) ;
    dffr camera_module_cache_reg_ram_233__5 (.Q (camera_module_cache_ram_233__5)
         , .QB (\$dummy [1724]), .D (nx15083), .CLK (clk), .R (rst)) ;
    mux21_ni ix15084 (.Y (nx15083), .A0 (camera_module_cache_ram_233__5), .A1 (
             nx35488), .S0 (nx34448)) ;
    dffr camera_module_cache_reg_ram_249__5 (.Q (camera_module_cache_ram_249__5)
         , .QB (\$dummy [1725]), .D (nx15073), .CLK (clk), .R (rst)) ;
    mux21_ni ix15074 (.Y (nx15073), .A0 (camera_module_cache_ram_249__5), .A1 (
             nx35488), .S0 (nx34444)) ;
    oai21 ix31832 (.Y (nx31831), .A0 (nx18168), .A1 (nx18090), .B0 (nx36488)) ;
    nand04 ix18169 (.Y (nx18168), .A0 (nx31834), .A1 (nx31842), .A2 (nx31850), .A3 (
           nx31858)) ;
    aoi22 ix31835 (.Y (nx31834), .A0 (camera_module_cache_ram_10__5), .A1 (
          nx35838), .B0 (camera_module_cache_ram_26__5), .B1 (nx35878)) ;
    dffr camera_module_cache_reg_ram_10__5 (.Q (camera_module_cache_ram_10__5), 
         .QB (\$dummy [1726]), .D (nx15063), .CLK (clk), .R (rst)) ;
    mux21_ni ix15064 (.Y (nx15063), .A0 (camera_module_cache_ram_10__5), .A1 (
             nx35488), .S0 (nx34434)) ;
    dffr camera_module_cache_reg_ram_26__5 (.Q (camera_module_cache_ram_26__5), 
         .QB (\$dummy [1727]), .D (nx15053), .CLK (clk), .R (rst)) ;
    mux21_ni ix15054 (.Y (nx15053), .A0 (camera_module_cache_ram_26__5), .A1 (
             nx35490), .S0 (nx34430)) ;
    aoi22 ix31843 (.Y (nx31842), .A0 (camera_module_cache_ram_42__5), .A1 (
          nx35918), .B0 (camera_module_cache_ram_58__5), .B1 (nx35958)) ;
    dffr camera_module_cache_reg_ram_42__5 (.Q (camera_module_cache_ram_42__5), 
         .QB (\$dummy [1728]), .D (nx15043), .CLK (clk), .R (rst)) ;
    mux21_ni ix15044 (.Y (nx15043), .A0 (camera_module_cache_ram_42__5), .A1 (
             nx35490), .S0 (nx34426)) ;
    dffr camera_module_cache_reg_ram_58__5 (.Q (camera_module_cache_ram_58__5), 
         .QB (\$dummy [1729]), .D (nx15033), .CLK (clk), .R (rst)) ;
    mux21_ni ix15034 (.Y (nx15033), .A0 (camera_module_cache_ram_58__5), .A1 (
             nx35490), .S0 (nx34422)) ;
    aoi22 ix31851 (.Y (nx31850), .A0 (camera_module_cache_ram_74__5), .A1 (
          nx35998), .B0 (camera_module_cache_ram_90__5), .B1 (nx36038)) ;
    dffr camera_module_cache_reg_ram_74__5 (.Q (camera_module_cache_ram_74__5), 
         .QB (\$dummy [1730]), .D (nx15023), .CLK (clk), .R (rst)) ;
    mux21_ni ix15024 (.Y (nx15023), .A0 (camera_module_cache_ram_74__5), .A1 (
             nx35490), .S0 (nx34418)) ;
    dffr camera_module_cache_reg_ram_90__5 (.Q (camera_module_cache_ram_90__5), 
         .QB (\$dummy [1731]), .D (nx15013), .CLK (clk), .R (rst)) ;
    mux21_ni ix15014 (.Y (nx15013), .A0 (camera_module_cache_ram_90__5), .A1 (
             nx35490), .S0 (nx34414)) ;
    aoi22 ix31859 (.Y (nx31858), .A0 (camera_module_cache_ram_122__5), .A1 (
          nx36078), .B0 (camera_module_cache_ram_106__5), .B1 (nx36118)) ;
    dffr camera_module_cache_reg_ram_122__5 (.Q (camera_module_cache_ram_122__5)
         , .QB (\$dummy [1732]), .D (nx14993), .CLK (clk), .R (rst)) ;
    mux21_ni ix14994 (.Y (nx14993), .A0 (camera_module_cache_ram_122__5), .A1 (
             nx35490), .S0 (nx34406)) ;
    dffr camera_module_cache_reg_ram_106__5 (.Q (camera_module_cache_ram_106__5)
         , .QB (\$dummy [1733]), .D (nx15003), .CLK (clk), .R (rst)) ;
    mux21_ni ix15004 (.Y (nx15003), .A0 (camera_module_cache_ram_106__5), .A1 (
             nx35490), .S0 (nx34410)) ;
    nand04 ix18091 (.Y (nx18090), .A0 (nx31867), .A1 (nx31875), .A2 (nx31883), .A3 (
           nx31891)) ;
    aoi22 ix31868 (.Y (nx31867), .A0 (camera_module_cache_ram_138__5), .A1 (
          nx36158), .B0 (camera_module_cache_ram_154__5), .B1 (nx36198)) ;
    dffr camera_module_cache_reg_ram_138__5 (.Q (camera_module_cache_ram_138__5)
         , .QB (\$dummy [1734]), .D (nx14983), .CLK (clk), .R (rst)) ;
    mux21_ni ix14984 (.Y (nx14983), .A0 (camera_module_cache_ram_138__5), .A1 (
             nx35492), .S0 (nx34402)) ;
    dffr camera_module_cache_reg_ram_154__5 (.Q (camera_module_cache_ram_154__5)
         , .QB (\$dummy [1735]), .D (nx14973), .CLK (clk), .R (rst)) ;
    mux21_ni ix14974 (.Y (nx14973), .A0 (camera_module_cache_ram_154__5), .A1 (
             nx35492), .S0 (nx34398)) ;
    aoi22 ix31876 (.Y (nx31875), .A0 (camera_module_cache_ram_186__5), .A1 (
          nx36238), .B0 (camera_module_cache_ram_170__5), .B1 (nx36278)) ;
    dffr camera_module_cache_reg_ram_186__5 (.Q (camera_module_cache_ram_186__5)
         , .QB (\$dummy [1736]), .D (nx14953), .CLK (clk), .R (rst)) ;
    mux21_ni ix14954 (.Y (nx14953), .A0 (camera_module_cache_ram_186__5), .A1 (
             nx35492), .S0 (nx34390)) ;
    dffr camera_module_cache_reg_ram_170__5 (.Q (camera_module_cache_ram_170__5)
         , .QB (\$dummy [1737]), .D (nx14963), .CLK (clk), .R (rst)) ;
    mux21_ni ix14964 (.Y (nx14963), .A0 (camera_module_cache_ram_170__5), .A1 (
             nx35492), .S0 (nx34394)) ;
    aoi22 ix31884 (.Y (nx31883), .A0 (camera_module_cache_ram_202__5), .A1 (
          nx36318), .B0 (camera_module_cache_ram_218__5), .B1 (nx36358)) ;
    dffr camera_module_cache_reg_ram_202__5 (.Q (camera_module_cache_ram_202__5)
         , .QB (\$dummy [1738]), .D (nx14943), .CLK (clk), .R (rst)) ;
    mux21_ni ix14944 (.Y (nx14943), .A0 (camera_module_cache_ram_202__5), .A1 (
             nx35492), .S0 (nx34386)) ;
    dffr camera_module_cache_reg_ram_218__5 (.Q (camera_module_cache_ram_218__5)
         , .QB (\$dummy [1739]), .D (nx14933), .CLK (clk), .R (rst)) ;
    mux21_ni ix14934 (.Y (nx14933), .A0 (camera_module_cache_ram_218__5), .A1 (
             nx35492), .S0 (nx34382)) ;
    aoi22 ix31892 (.Y (nx31891), .A0 (camera_module_cache_ram_234__5), .A1 (
          nx36398), .B0 (camera_module_cache_ram_250__5), .B1 (nx36438)) ;
    dffr camera_module_cache_reg_ram_234__5 (.Q (camera_module_cache_ram_234__5)
         , .QB (\$dummy [1740]), .D (nx14923), .CLK (clk), .R (rst)) ;
    mux21_ni ix14924 (.Y (nx14923), .A0 (camera_module_cache_ram_234__5), .A1 (
             nx35492), .S0 (nx34378)) ;
    dffr camera_module_cache_reg_ram_250__5 (.Q (camera_module_cache_ram_250__5)
         , .QB (\$dummy [1741]), .D (nx14913), .CLK (clk), .R (rst)) ;
    mux21_ni ix14914 (.Y (nx14913), .A0 (camera_module_cache_ram_250__5), .A1 (
             nx35494), .S0 (nx34374)) ;
    oai21 ix31900 (.Y (nx31899), .A0 (nx18006), .A1 (nx17928), .B0 (nx36492)) ;
    nand04 ix18007 (.Y (nx18006), .A0 (nx31902), .A1 (nx31910), .A2 (nx31918), .A3 (
           nx31926)) ;
    aoi22 ix31903 (.Y (nx31902), .A0 (camera_module_cache_ram_11__5), .A1 (
          nx35838), .B0 (camera_module_cache_ram_27__5), .B1 (nx35878)) ;
    dffr camera_module_cache_reg_ram_11__5 (.Q (camera_module_cache_ram_11__5), 
         .QB (\$dummy [1742]), .D (nx14903), .CLK (clk), .R (rst)) ;
    mux21_ni ix14904 (.Y (nx14903), .A0 (camera_module_cache_ram_11__5), .A1 (
             nx35494), .S0 (nx34364)) ;
    dffr camera_module_cache_reg_ram_27__5 (.Q (camera_module_cache_ram_27__5), 
         .QB (\$dummy [1743]), .D (nx14893), .CLK (clk), .R (rst)) ;
    mux21_ni ix14894 (.Y (nx14893), .A0 (camera_module_cache_ram_27__5), .A1 (
             nx35494), .S0 (nx34360)) ;
    aoi22 ix31911 (.Y (nx31910), .A0 (camera_module_cache_ram_43__5), .A1 (
          nx35918), .B0 (camera_module_cache_ram_59__5), .B1 (nx35958)) ;
    dffr camera_module_cache_reg_ram_43__5 (.Q (camera_module_cache_ram_43__5), 
         .QB (\$dummy [1744]), .D (nx14883), .CLK (clk), .R (rst)) ;
    mux21_ni ix14884 (.Y (nx14883), .A0 (camera_module_cache_ram_43__5), .A1 (
             nx35494), .S0 (nx34356)) ;
    dffr camera_module_cache_reg_ram_59__5 (.Q (camera_module_cache_ram_59__5), 
         .QB (\$dummy [1745]), .D (nx14873), .CLK (clk), .R (rst)) ;
    mux21_ni ix14874 (.Y (nx14873), .A0 (camera_module_cache_ram_59__5), .A1 (
             nx35494), .S0 (nx34352)) ;
    aoi22 ix31919 (.Y (nx31918), .A0 (camera_module_cache_ram_75__5), .A1 (
          nx35998), .B0 (camera_module_cache_ram_91__5), .B1 (nx36038)) ;
    dffr camera_module_cache_reg_ram_75__5 (.Q (camera_module_cache_ram_75__5), 
         .QB (\$dummy [1746]), .D (nx14863), .CLK (clk), .R (rst)) ;
    mux21_ni ix14864 (.Y (nx14863), .A0 (camera_module_cache_ram_75__5), .A1 (
             nx35494), .S0 (nx34348)) ;
    dffr camera_module_cache_reg_ram_91__5 (.Q (camera_module_cache_ram_91__5), 
         .QB (\$dummy [1747]), .D (nx14853), .CLK (clk), .R (rst)) ;
    mux21_ni ix14854 (.Y (nx14853), .A0 (camera_module_cache_ram_91__5), .A1 (
             nx35494), .S0 (nx34344)) ;
    aoi22 ix31927 (.Y (nx31926), .A0 (camera_module_cache_ram_123__5), .A1 (
          nx36078), .B0 (camera_module_cache_ram_107__5), .B1 (nx36118)) ;
    dffr camera_module_cache_reg_ram_123__5 (.Q (camera_module_cache_ram_123__5)
         , .QB (\$dummy [1748]), .D (nx14833), .CLK (clk), .R (rst)) ;
    mux21_ni ix14834 (.Y (nx14833), .A0 (camera_module_cache_ram_123__5), .A1 (
             nx35496), .S0 (nx34336)) ;
    dffr camera_module_cache_reg_ram_107__5 (.Q (camera_module_cache_ram_107__5)
         , .QB (\$dummy [1749]), .D (nx14843), .CLK (clk), .R (rst)) ;
    mux21_ni ix14844 (.Y (nx14843), .A0 (camera_module_cache_ram_107__5), .A1 (
             nx35496), .S0 (nx34340)) ;
    nand04 ix17929 (.Y (nx17928), .A0 (nx31935), .A1 (nx31943), .A2 (nx31951), .A3 (
           nx31959)) ;
    aoi22 ix31936 (.Y (nx31935), .A0 (camera_module_cache_ram_139__5), .A1 (
          nx36158), .B0 (camera_module_cache_ram_155__5), .B1 (nx36198)) ;
    dffr camera_module_cache_reg_ram_139__5 (.Q (camera_module_cache_ram_139__5)
         , .QB (\$dummy [1750]), .D (nx14823), .CLK (clk), .R (rst)) ;
    mux21_ni ix14824 (.Y (nx14823), .A0 (camera_module_cache_ram_139__5), .A1 (
             nx35496), .S0 (nx34332)) ;
    dffr camera_module_cache_reg_ram_155__5 (.Q (camera_module_cache_ram_155__5)
         , .QB (\$dummy [1751]), .D (nx14813), .CLK (clk), .R (rst)) ;
    mux21_ni ix14814 (.Y (nx14813), .A0 (camera_module_cache_ram_155__5), .A1 (
             nx35496), .S0 (nx34328)) ;
    aoi22 ix31944 (.Y (nx31943), .A0 (camera_module_cache_ram_187__5), .A1 (
          nx36238), .B0 (camera_module_cache_ram_171__5), .B1 (nx36278)) ;
    dffr camera_module_cache_reg_ram_187__5 (.Q (camera_module_cache_ram_187__5)
         , .QB (\$dummy [1752]), .D (nx14793), .CLK (clk), .R (rst)) ;
    mux21_ni ix14794 (.Y (nx14793), .A0 (camera_module_cache_ram_187__5), .A1 (
             nx35496), .S0 (nx34320)) ;
    dffr camera_module_cache_reg_ram_171__5 (.Q (camera_module_cache_ram_171__5)
         , .QB (\$dummy [1753]), .D (nx14803), .CLK (clk), .R (rst)) ;
    mux21_ni ix14804 (.Y (nx14803), .A0 (camera_module_cache_ram_171__5), .A1 (
             nx35496), .S0 (nx34324)) ;
    aoi22 ix31952 (.Y (nx31951), .A0 (camera_module_cache_ram_203__5), .A1 (
          nx36318), .B0 (camera_module_cache_ram_219__5), .B1 (nx36358)) ;
    dffr camera_module_cache_reg_ram_203__5 (.Q (camera_module_cache_ram_203__5)
         , .QB (\$dummy [1754]), .D (nx14783), .CLK (clk), .R (rst)) ;
    mux21_ni ix14784 (.Y (nx14783), .A0 (camera_module_cache_ram_203__5), .A1 (
             nx35496), .S0 (nx34316)) ;
    dffr camera_module_cache_reg_ram_219__5 (.Q (camera_module_cache_ram_219__5)
         , .QB (\$dummy [1755]), .D (nx14773), .CLK (clk), .R (rst)) ;
    mux21_ni ix14774 (.Y (nx14773), .A0 (camera_module_cache_ram_219__5), .A1 (
             nx35498), .S0 (nx34312)) ;
    aoi22 ix31960 (.Y (nx31959), .A0 (camera_module_cache_ram_235__5), .A1 (
          nx36398), .B0 (camera_module_cache_ram_251__5), .B1 (nx36438)) ;
    dffr camera_module_cache_reg_ram_235__5 (.Q (camera_module_cache_ram_235__5)
         , .QB (\$dummy [1756]), .D (nx14763), .CLK (clk), .R (rst)) ;
    mux21_ni ix14764 (.Y (nx14763), .A0 (camera_module_cache_ram_235__5), .A1 (
             nx35498), .S0 (nx34308)) ;
    dffr camera_module_cache_reg_ram_251__5 (.Q (camera_module_cache_ram_251__5)
         , .QB (\$dummy [1757]), .D (nx14753), .CLK (clk), .R (rst)) ;
    mux21_ni ix14754 (.Y (nx14753), .A0 (camera_module_cache_ram_251__5), .A1 (
             nx35498), .S0 (nx34304)) ;
    nand04 ix17851 (.Y (nx17850), .A0 (nx31968), .A1 (nx32036), .A2 (nx32104), .A3 (
           nx32172)) ;
    oai21 ix31969 (.Y (nx31968), .A0 (nx17840), .A1 (nx17762), .B0 (nx36508)) ;
    nand04 ix17841 (.Y (nx17840), .A0 (nx31971), .A1 (nx31979), .A2 (nx31987), .A3 (
           nx31995)) ;
    aoi22 ix31972 (.Y (nx31971), .A0 (camera_module_cache_ram_12__5), .A1 (
          nx35840), .B0 (camera_module_cache_ram_28__5), .B1 (nx35880)) ;
    dffr camera_module_cache_reg_ram_12__5 (.Q (camera_module_cache_ram_12__5), 
         .QB (\$dummy [1758]), .D (nx14743), .CLK (clk), .R (rst)) ;
    mux21_ni ix14744 (.Y (nx14743), .A0 (nx35498), .A1 (
             camera_module_cache_ram_12__5), .S0 (nx36496)) ;
    dffr camera_module_cache_reg_ram_28__5 (.Q (camera_module_cache_ram_28__5), 
         .QB (\$dummy [1759]), .D (nx14733), .CLK (clk), .R (rst)) ;
    mux21_ni ix14734 (.Y (nx14733), .A0 (nx35498), .A1 (
             camera_module_cache_ram_28__5), .S0 (nx36510)) ;
    aoi22 ix31980 (.Y (nx31979), .A0 (camera_module_cache_ram_44__5), .A1 (
          nx35920), .B0 (camera_module_cache_ram_60__5), .B1 (nx35960)) ;
    dffr camera_module_cache_reg_ram_44__5 (.Q (camera_module_cache_ram_44__5), 
         .QB (\$dummy [1760]), .D (nx14723), .CLK (clk), .R (rst)) ;
    mux21_ni ix14724 (.Y (nx14723), .A0 (nx35498), .A1 (
             camera_module_cache_ram_44__5), .S0 (nx36514)) ;
    dffr camera_module_cache_reg_ram_60__5 (.Q (camera_module_cache_ram_60__5), 
         .QB (\$dummy [1761]), .D (nx14713), .CLK (clk), .R (rst)) ;
    mux21_ni ix14714 (.Y (nx14713), .A0 (nx35498), .A1 (
             camera_module_cache_ram_60__5), .S0 (nx36518)) ;
    aoi22 ix31988 (.Y (nx31987), .A0 (camera_module_cache_ram_76__5), .A1 (
          nx36000), .B0 (camera_module_cache_ram_92__5), .B1 (nx36040)) ;
    dffr camera_module_cache_reg_ram_76__5 (.Q (camera_module_cache_ram_76__5), 
         .QB (\$dummy [1762]), .D (nx14703), .CLK (clk), .R (rst)) ;
    mux21_ni ix14704 (.Y (nx14703), .A0 (nx35500), .A1 (
             camera_module_cache_ram_76__5), .S0 (nx36522)) ;
    dffr camera_module_cache_reg_ram_92__5 (.Q (camera_module_cache_ram_92__5), 
         .QB (\$dummy [1763]), .D (nx14693), .CLK (clk), .R (rst)) ;
    mux21_ni ix14694 (.Y (nx14693), .A0 (nx35500), .A1 (
             camera_module_cache_ram_92__5), .S0 (nx36526)) ;
    aoi22 ix31996 (.Y (nx31995), .A0 (camera_module_cache_ram_124__5), .A1 (
          nx36080), .B0 (camera_module_cache_ram_108__5), .B1 (nx36120)) ;
    dffr camera_module_cache_reg_ram_124__5 (.Q (camera_module_cache_ram_124__5)
         , .QB (\$dummy [1764]), .D (nx14673), .CLK (clk), .R (rst)) ;
    mux21_ni ix14674 (.Y (nx14673), .A0 (nx35500), .A1 (
             camera_module_cache_ram_124__5), .S0 (nx36530)) ;
    dffr camera_module_cache_reg_ram_108__5 (.Q (camera_module_cache_ram_108__5)
         , .QB (\$dummy [1765]), .D (nx14683), .CLK (clk), .R (rst)) ;
    mux21_ni ix14684 (.Y (nx14683), .A0 (nx35500), .A1 (
             camera_module_cache_ram_108__5), .S0 (nx36534)) ;
    nand04 ix17763 (.Y (nx17762), .A0 (nx32004), .A1 (nx32012), .A2 (nx32020), .A3 (
           nx32028)) ;
    aoi22 ix32005 (.Y (nx32004), .A0 (camera_module_cache_ram_140__5), .A1 (
          nx36160), .B0 (camera_module_cache_ram_156__5), .B1 (nx36200)) ;
    dffr camera_module_cache_reg_ram_140__5 (.Q (camera_module_cache_ram_140__5)
         , .QB (\$dummy [1766]), .D (nx14663), .CLK (clk), .R (rst)) ;
    mux21_ni ix14664 (.Y (nx14663), .A0 (nx35500), .A1 (
             camera_module_cache_ram_140__5), .S0 (nx36538)) ;
    dffr camera_module_cache_reg_ram_156__5 (.Q (camera_module_cache_ram_156__5)
         , .QB (\$dummy [1767]), .D (nx14653), .CLK (clk), .R (rst)) ;
    mux21_ni ix14654 (.Y (nx14653), .A0 (nx35500), .A1 (
             camera_module_cache_ram_156__5), .S0 (nx36542)) ;
    aoi22 ix32013 (.Y (nx32012), .A0 (camera_module_cache_ram_188__5), .A1 (
          nx36240), .B0 (camera_module_cache_ram_172__5), .B1 (nx36280)) ;
    dffr camera_module_cache_reg_ram_188__5 (.Q (camera_module_cache_ram_188__5)
         , .QB (\$dummy [1768]), .D (nx14633), .CLK (clk), .R (rst)) ;
    mux21_ni ix14634 (.Y (nx14633), .A0 (nx35500), .A1 (
             camera_module_cache_ram_188__5), .S0 (nx36546)) ;
    dffr camera_module_cache_reg_ram_172__5 (.Q (camera_module_cache_ram_172__5)
         , .QB (\$dummy [1769]), .D (nx14643), .CLK (clk), .R (rst)) ;
    mux21_ni ix14644 (.Y (nx14643), .A0 (nx35502), .A1 (
             camera_module_cache_ram_172__5), .S0 (nx36550)) ;
    aoi22 ix32021 (.Y (nx32020), .A0 (camera_module_cache_ram_204__5), .A1 (
          nx36320), .B0 (camera_module_cache_ram_220__5), .B1 (nx36360)) ;
    dffr camera_module_cache_reg_ram_204__5 (.Q (camera_module_cache_ram_204__5)
         , .QB (\$dummy [1770]), .D (nx14623), .CLK (clk), .R (rst)) ;
    mux21_ni ix14624 (.Y (nx14623), .A0 (nx35502), .A1 (
             camera_module_cache_ram_204__5), .S0 (nx36554)) ;
    dffr camera_module_cache_reg_ram_220__5 (.Q (camera_module_cache_ram_220__5)
         , .QB (\$dummy [1771]), .D (nx14613), .CLK (clk), .R (rst)) ;
    mux21_ni ix14614 (.Y (nx14613), .A0 (nx35502), .A1 (
             camera_module_cache_ram_220__5), .S0 (nx36558)) ;
    aoi22 ix32029 (.Y (nx32028), .A0 (camera_module_cache_ram_236__5), .A1 (
          nx36400), .B0 (camera_module_cache_ram_252__5), .B1 (nx36440)) ;
    dffr camera_module_cache_reg_ram_236__5 (.Q (camera_module_cache_ram_236__5)
         , .QB (\$dummy [1772]), .D (nx14603), .CLK (clk), .R (rst)) ;
    mux21_ni ix14604 (.Y (nx14603), .A0 (nx35502), .A1 (
             camera_module_cache_ram_236__5), .S0 (nx36562)) ;
    dffr camera_module_cache_reg_ram_252__5 (.Q (camera_module_cache_ram_252__5)
         , .QB (\$dummy [1773]), .D (nx14593), .CLK (clk), .R (rst)) ;
    mux21_ni ix14594 (.Y (nx14593), .A0 (nx35502), .A1 (
             camera_module_cache_ram_252__5), .S0 (nx36566)) ;
    oai21 ix32037 (.Y (nx32036), .A0 (nx17678), .A1 (nx17600), .B0 (nx36582)) ;
    nand04 ix17679 (.Y (nx17678), .A0 (nx32039), .A1 (nx32047), .A2 (nx32055), .A3 (
           nx32063)) ;
    aoi22 ix32040 (.Y (nx32039), .A0 (camera_module_cache_ram_13__5), .A1 (
          nx35840), .B0 (camera_module_cache_ram_29__5), .B1 (nx35880)) ;
    dffr camera_module_cache_reg_ram_13__5 (.Q (camera_module_cache_ram_13__5), 
         .QB (\$dummy [1774]), .D (nx14583), .CLK (clk), .R (rst)) ;
    mux21_ni ix14584 (.Y (nx14583), .A0 (nx35502), .A1 (
             camera_module_cache_ram_13__5), .S0 (nx36570)) ;
    dffr camera_module_cache_reg_ram_29__5 (.Q (camera_module_cache_ram_29__5), 
         .QB (\$dummy [1775]), .D (nx14573), .CLK (clk), .R (rst)) ;
    mux21_ni ix14574 (.Y (nx14573), .A0 (nx35502), .A1 (
             camera_module_cache_ram_29__5), .S0 (nx36584)) ;
    aoi22 ix32048 (.Y (nx32047), .A0 (camera_module_cache_ram_45__5), .A1 (
          nx35920), .B0 (camera_module_cache_ram_61__5), .B1 (nx35960)) ;
    dffr camera_module_cache_reg_ram_45__5 (.Q (camera_module_cache_ram_45__5), 
         .QB (\$dummy [1776]), .D (nx14563), .CLK (clk), .R (rst)) ;
    mux21_ni ix14564 (.Y (nx14563), .A0 (nx35504), .A1 (
             camera_module_cache_ram_45__5), .S0 (nx36588)) ;
    dffr camera_module_cache_reg_ram_61__5 (.Q (camera_module_cache_ram_61__5), 
         .QB (\$dummy [1777]), .D (nx14553), .CLK (clk), .R (rst)) ;
    mux21_ni ix14554 (.Y (nx14553), .A0 (nx35504), .A1 (
             camera_module_cache_ram_61__5), .S0 (nx36592)) ;
    aoi22 ix32056 (.Y (nx32055), .A0 (camera_module_cache_ram_77__5), .A1 (
          nx36000), .B0 (camera_module_cache_ram_93__5), .B1 (nx36040)) ;
    dffr camera_module_cache_reg_ram_77__5 (.Q (camera_module_cache_ram_77__5), 
         .QB (\$dummy [1778]), .D (nx14543), .CLK (clk), .R (rst)) ;
    mux21_ni ix14544 (.Y (nx14543), .A0 (nx35504), .A1 (
             camera_module_cache_ram_77__5), .S0 (nx36596)) ;
    dffr camera_module_cache_reg_ram_93__5 (.Q (camera_module_cache_ram_93__5), 
         .QB (\$dummy [1779]), .D (nx14533), .CLK (clk), .R (rst)) ;
    mux21_ni ix14534 (.Y (nx14533), .A0 (nx35504), .A1 (
             camera_module_cache_ram_93__5), .S0 (nx36600)) ;
    aoi22 ix32064 (.Y (nx32063), .A0 (camera_module_cache_ram_125__5), .A1 (
          nx36080), .B0 (camera_module_cache_ram_109__5), .B1 (nx36120)) ;
    dffr camera_module_cache_reg_ram_125__5 (.Q (camera_module_cache_ram_125__5)
         , .QB (\$dummy [1780]), .D (nx14513), .CLK (clk), .R (rst)) ;
    mux21_ni ix14514 (.Y (nx14513), .A0 (nx35504), .A1 (
             camera_module_cache_ram_125__5), .S0 (nx36604)) ;
    dffr camera_module_cache_reg_ram_109__5 (.Q (camera_module_cache_ram_109__5)
         , .QB (\$dummy [1781]), .D (nx14523), .CLK (clk), .R (rst)) ;
    mux21_ni ix14524 (.Y (nx14523), .A0 (nx35504), .A1 (
             camera_module_cache_ram_109__5), .S0 (nx36608)) ;
    nand04 ix17601 (.Y (nx17600), .A0 (nx32072), .A1 (nx32080), .A2 (nx32088), .A3 (
           nx32096)) ;
    aoi22 ix32073 (.Y (nx32072), .A0 (camera_module_cache_ram_141__5), .A1 (
          nx36160), .B0 (camera_module_cache_ram_157__5), .B1 (nx36200)) ;
    dffr camera_module_cache_reg_ram_141__5 (.Q (camera_module_cache_ram_141__5)
         , .QB (\$dummy [1782]), .D (nx14503), .CLK (clk), .R (rst)) ;
    mux21_ni ix14504 (.Y (nx14503), .A0 (nx35504), .A1 (
             camera_module_cache_ram_141__5), .S0 (nx36612)) ;
    dffr camera_module_cache_reg_ram_157__5 (.Q (camera_module_cache_ram_157__5)
         , .QB (\$dummy [1783]), .D (nx14493), .CLK (clk), .R (rst)) ;
    mux21_ni ix14494 (.Y (nx14493), .A0 (nx35506), .A1 (
             camera_module_cache_ram_157__5), .S0 (nx36616)) ;
    aoi22 ix32081 (.Y (nx32080), .A0 (camera_module_cache_ram_189__5), .A1 (
          nx36240), .B0 (camera_module_cache_ram_173__5), .B1 (nx36280)) ;
    dffr camera_module_cache_reg_ram_189__5 (.Q (camera_module_cache_ram_189__5)
         , .QB (\$dummy [1784]), .D (nx14473), .CLK (clk), .R (rst)) ;
    mux21_ni ix14474 (.Y (nx14473), .A0 (nx35506), .A1 (
             camera_module_cache_ram_189__5), .S0 (nx36620)) ;
    dffr camera_module_cache_reg_ram_173__5 (.Q (camera_module_cache_ram_173__5)
         , .QB (\$dummy [1785]), .D (nx14483), .CLK (clk), .R (rst)) ;
    mux21_ni ix14484 (.Y (nx14483), .A0 (nx35506), .A1 (
             camera_module_cache_ram_173__5), .S0 (nx36624)) ;
    aoi22 ix32089 (.Y (nx32088), .A0 (camera_module_cache_ram_205__5), .A1 (
          nx36320), .B0 (camera_module_cache_ram_221__5), .B1 (nx36360)) ;
    dffr camera_module_cache_reg_ram_205__5 (.Q (camera_module_cache_ram_205__5)
         , .QB (\$dummy [1786]), .D (nx14463), .CLK (clk), .R (rst)) ;
    mux21_ni ix14464 (.Y (nx14463), .A0 (nx35506), .A1 (
             camera_module_cache_ram_205__5), .S0 (nx36628)) ;
    dffr camera_module_cache_reg_ram_221__5 (.Q (camera_module_cache_ram_221__5)
         , .QB (\$dummy [1787]), .D (nx14453), .CLK (clk), .R (rst)) ;
    mux21_ni ix14454 (.Y (nx14453), .A0 (nx35506), .A1 (
             camera_module_cache_ram_221__5), .S0 (nx36632)) ;
    aoi22 ix32097 (.Y (nx32096), .A0 (camera_module_cache_ram_237__5), .A1 (
          nx36400), .B0 (camera_module_cache_ram_253__5), .B1 (nx36440)) ;
    dffr camera_module_cache_reg_ram_237__5 (.Q (camera_module_cache_ram_237__5)
         , .QB (\$dummy [1788]), .D (nx14443), .CLK (clk), .R (rst)) ;
    mux21_ni ix14444 (.Y (nx14443), .A0 (nx35506), .A1 (
             camera_module_cache_ram_237__5), .S0 (nx36636)) ;
    dffr camera_module_cache_reg_ram_253__5 (.Q (camera_module_cache_ram_253__5)
         , .QB (\$dummy [1789]), .D (nx14433), .CLK (clk), .R (rst)) ;
    mux21_ni ix14434 (.Y (nx14433), .A0 (nx35506), .A1 (
             camera_module_cache_ram_253__5), .S0 (nx36640)) ;
    oai21 ix32105 (.Y (nx32104), .A0 (nx17514), .A1 (nx17436), .B0 (nx36656)) ;
    nand04 ix17515 (.Y (nx17514), .A0 (nx32107), .A1 (nx32115), .A2 (nx32123), .A3 (
           nx32131)) ;
    aoi22 ix32108 (.Y (nx32107), .A0 (camera_module_cache_ram_14__5), .A1 (
          nx35840), .B0 (camera_module_cache_ram_30__5), .B1 (nx35880)) ;
    dffr camera_module_cache_reg_ram_14__5 (.Q (camera_module_cache_ram_14__5), 
         .QB (\$dummy [1790]), .D (nx14423), .CLK (clk), .R (rst)) ;
    mux21_ni ix14424 (.Y (nx14423), .A0 (nx35508), .A1 (
             camera_module_cache_ram_14__5), .S0 (nx36644)) ;
    dffr camera_module_cache_reg_ram_30__5 (.Q (camera_module_cache_ram_30__5), 
         .QB (\$dummy [1791]), .D (nx14413), .CLK (clk), .R (rst)) ;
    mux21_ni ix14414 (.Y (nx14413), .A0 (nx35508), .A1 (
             camera_module_cache_ram_30__5), .S0 (nx36658)) ;
    aoi22 ix32116 (.Y (nx32115), .A0 (camera_module_cache_ram_46__5), .A1 (
          nx35920), .B0 (camera_module_cache_ram_62__5), .B1 (nx35960)) ;
    dffr camera_module_cache_reg_ram_46__5 (.Q (camera_module_cache_ram_46__5), 
         .QB (\$dummy [1792]), .D (nx14403), .CLK (clk), .R (rst)) ;
    mux21_ni ix14404 (.Y (nx14403), .A0 (nx35508), .A1 (
             camera_module_cache_ram_46__5), .S0 (nx36662)) ;
    dffr camera_module_cache_reg_ram_62__5 (.Q (camera_module_cache_ram_62__5), 
         .QB (\$dummy [1793]), .D (nx14393), .CLK (clk), .R (rst)) ;
    mux21_ni ix14394 (.Y (nx14393), .A0 (nx35508), .A1 (
             camera_module_cache_ram_62__5), .S0 (nx36666)) ;
    aoi22 ix32124 (.Y (nx32123), .A0 (camera_module_cache_ram_78__5), .A1 (
          nx36000), .B0 (camera_module_cache_ram_94__5), .B1 (nx36040)) ;
    dffr camera_module_cache_reg_ram_78__5 (.Q (camera_module_cache_ram_78__5), 
         .QB (\$dummy [1794]), .D (nx14383), .CLK (clk), .R (rst)) ;
    mux21_ni ix14384 (.Y (nx14383), .A0 (nx35508), .A1 (
             camera_module_cache_ram_78__5), .S0 (nx36670)) ;
    dffr camera_module_cache_reg_ram_94__5 (.Q (camera_module_cache_ram_94__5), 
         .QB (\$dummy [1795]), .D (nx14373), .CLK (clk), .R (rst)) ;
    mux21_ni ix14374 (.Y (nx14373), .A0 (nx35508), .A1 (
             camera_module_cache_ram_94__5), .S0 (nx36674)) ;
    aoi22 ix32132 (.Y (nx32131), .A0 (camera_module_cache_ram_126__5), .A1 (
          nx36080), .B0 (camera_module_cache_ram_110__5), .B1 (nx36120)) ;
    dffr camera_module_cache_reg_ram_126__5 (.Q (camera_module_cache_ram_126__5)
         , .QB (\$dummy [1796]), .D (nx14353), .CLK (clk), .R (rst)) ;
    mux21_ni ix14354 (.Y (nx14353), .A0 (nx35508), .A1 (
             camera_module_cache_ram_126__5), .S0 (nx36678)) ;
    dffr camera_module_cache_reg_ram_110__5 (.Q (camera_module_cache_ram_110__5)
         , .QB (\$dummy [1797]), .D (nx14363), .CLK (clk), .R (rst)) ;
    mux21_ni ix14364 (.Y (nx14363), .A0 (nx35510), .A1 (
             camera_module_cache_ram_110__5), .S0 (nx36682)) ;
    nand04 ix17437 (.Y (nx17436), .A0 (nx32140), .A1 (nx32148), .A2 (nx32156), .A3 (
           nx32164)) ;
    aoi22 ix32141 (.Y (nx32140), .A0 (camera_module_cache_ram_142__5), .A1 (
          nx36160), .B0 (camera_module_cache_ram_158__5), .B1 (nx36200)) ;
    dffr camera_module_cache_reg_ram_142__5 (.Q (camera_module_cache_ram_142__5)
         , .QB (\$dummy [1798]), .D (nx14343), .CLK (clk), .R (rst)) ;
    mux21_ni ix14344 (.Y (nx14343), .A0 (nx35510), .A1 (
             camera_module_cache_ram_142__5), .S0 (nx36686)) ;
    dffr camera_module_cache_reg_ram_158__5 (.Q (camera_module_cache_ram_158__5)
         , .QB (\$dummy [1799]), .D (nx14333), .CLK (clk), .R (rst)) ;
    mux21_ni ix14334 (.Y (nx14333), .A0 (nx35510), .A1 (
             camera_module_cache_ram_158__5), .S0 (nx36690)) ;
    aoi22 ix32149 (.Y (nx32148), .A0 (camera_module_cache_ram_190__5), .A1 (
          nx36240), .B0 (camera_module_cache_ram_174__5), .B1 (nx36280)) ;
    dffr camera_module_cache_reg_ram_190__5 (.Q (camera_module_cache_ram_190__5)
         , .QB (\$dummy [1800]), .D (nx14313), .CLK (clk), .R (rst)) ;
    mux21_ni ix14314 (.Y (nx14313), .A0 (nx35510), .A1 (
             camera_module_cache_ram_190__5), .S0 (nx36694)) ;
    dffr camera_module_cache_reg_ram_174__5 (.Q (camera_module_cache_ram_174__5)
         , .QB (\$dummy [1801]), .D (nx14323), .CLK (clk), .R (rst)) ;
    mux21_ni ix14324 (.Y (nx14323), .A0 (nx35510), .A1 (
             camera_module_cache_ram_174__5), .S0 (nx36698)) ;
    aoi22 ix32157 (.Y (nx32156), .A0 (camera_module_cache_ram_206__5), .A1 (
          nx36320), .B0 (camera_module_cache_ram_222__5), .B1 (nx36360)) ;
    dffr camera_module_cache_reg_ram_206__5 (.Q (camera_module_cache_ram_206__5)
         , .QB (\$dummy [1802]), .D (nx14303), .CLK (clk), .R (rst)) ;
    mux21_ni ix14304 (.Y (nx14303), .A0 (nx35510), .A1 (
             camera_module_cache_ram_206__5), .S0 (nx36702)) ;
    dffr camera_module_cache_reg_ram_222__5 (.Q (camera_module_cache_ram_222__5)
         , .QB (\$dummy [1803]), .D (nx14293), .CLK (clk), .R (rst)) ;
    mux21_ni ix14294 (.Y (nx14293), .A0 (nx35510), .A1 (
             camera_module_cache_ram_222__5), .S0 (nx36706)) ;
    aoi22 ix32165 (.Y (nx32164), .A0 (camera_module_cache_ram_238__5), .A1 (
          nx36400), .B0 (camera_module_cache_ram_254__5), .B1 (nx36440)) ;
    dffr camera_module_cache_reg_ram_238__5 (.Q (camera_module_cache_ram_238__5)
         , .QB (\$dummy [1804]), .D (nx14283), .CLK (clk), .R (rst)) ;
    mux21_ni ix14284 (.Y (nx14283), .A0 (nx35512), .A1 (
             camera_module_cache_ram_238__5), .S0 (nx36710)) ;
    dffr camera_module_cache_reg_ram_254__5 (.Q (camera_module_cache_ram_254__5)
         , .QB (\$dummy [1805]), .D (nx14273), .CLK (clk), .R (rst)) ;
    mux21_ni ix14274 (.Y (nx14273), .A0 (nx35512), .A1 (
             camera_module_cache_ram_254__5), .S0 (nx36714)) ;
    oai21 ix32173 (.Y (nx32172), .A0 (nx17352), .A1 (nx17274), .B0 (nx36730)) ;
    nand04 ix17353 (.Y (nx17352), .A0 (nx32175), .A1 (nx32183), .A2 (nx32191), .A3 (
           nx32199)) ;
    aoi22 ix32176 (.Y (nx32175), .A0 (camera_module_cache_ram_15__5), .A1 (
          nx35840), .B0 (camera_module_cache_ram_31__5), .B1 (nx35880)) ;
    dffr camera_module_cache_reg_ram_15__5 (.Q (camera_module_cache_ram_15__5), 
         .QB (\$dummy [1806]), .D (nx14263), .CLK (clk), .R (rst)) ;
    mux21_ni ix14264 (.Y (nx14263), .A0 (nx35512), .A1 (
             camera_module_cache_ram_15__5), .S0 (nx36718)) ;
    dffr camera_module_cache_reg_ram_31__5 (.Q (camera_module_cache_ram_31__5), 
         .QB (\$dummy [1807]), .D (nx14253), .CLK (clk), .R (rst)) ;
    mux21_ni ix14254 (.Y (nx14253), .A0 (nx35512), .A1 (
             camera_module_cache_ram_31__5), .S0 (nx36732)) ;
    aoi22 ix32184 (.Y (nx32183), .A0 (camera_module_cache_ram_47__5), .A1 (
          nx35920), .B0 (camera_module_cache_ram_63__5), .B1 (nx35960)) ;
    dffr camera_module_cache_reg_ram_47__5 (.Q (camera_module_cache_ram_47__5), 
         .QB (\$dummy [1808]), .D (nx14243), .CLK (clk), .R (rst)) ;
    mux21_ni ix14244 (.Y (nx14243), .A0 (nx35512), .A1 (
             camera_module_cache_ram_47__5), .S0 (nx36736)) ;
    dffr camera_module_cache_reg_ram_63__5 (.Q (camera_module_cache_ram_63__5), 
         .QB (\$dummy [1809]), .D (nx14233), .CLK (clk), .R (rst)) ;
    mux21_ni ix14234 (.Y (nx14233), .A0 (nx35512), .A1 (
             camera_module_cache_ram_63__5), .S0 (nx36740)) ;
    aoi22 ix32192 (.Y (nx32191), .A0 (camera_module_cache_ram_79__5), .A1 (
          nx36000), .B0 (camera_module_cache_ram_95__5), .B1 (nx36040)) ;
    dffr camera_module_cache_reg_ram_79__5 (.Q (camera_module_cache_ram_79__5), 
         .QB (\$dummy [1810]), .D (nx14223), .CLK (clk), .R (rst)) ;
    mux21_ni ix14224 (.Y (nx14223), .A0 (nx35512), .A1 (
             camera_module_cache_ram_79__5), .S0 (nx36744)) ;
    dffr camera_module_cache_reg_ram_95__5 (.Q (camera_module_cache_ram_95__5), 
         .QB (\$dummy [1811]), .D (nx14213), .CLK (clk), .R (rst)) ;
    mux21_ni ix14214 (.Y (nx14213), .A0 (nx35514), .A1 (
             camera_module_cache_ram_95__5), .S0 (nx36748)) ;
    aoi22 ix32200 (.Y (nx32199), .A0 (camera_module_cache_ram_127__5), .A1 (
          nx36080), .B0 (camera_module_cache_ram_111__5), .B1 (nx36120)) ;
    dffr camera_module_cache_reg_ram_127__5 (.Q (camera_module_cache_ram_127__5)
         , .QB (\$dummy [1812]), .D (nx14193), .CLK (clk), .R (rst)) ;
    mux21_ni ix14194 (.Y (nx14193), .A0 (nx35514), .A1 (
             camera_module_cache_ram_127__5), .S0 (nx36752)) ;
    dffr camera_module_cache_reg_ram_111__5 (.Q (camera_module_cache_ram_111__5)
         , .QB (\$dummy [1813]), .D (nx14203), .CLK (clk), .R (rst)) ;
    mux21_ni ix14204 (.Y (nx14203), .A0 (nx35514), .A1 (
             camera_module_cache_ram_111__5), .S0 (nx36756)) ;
    nand04 ix17275 (.Y (nx17274), .A0 (nx32208), .A1 (nx32216), .A2 (nx32224), .A3 (
           nx32232)) ;
    aoi22 ix32209 (.Y (nx32208), .A0 (camera_module_cache_ram_143__5), .A1 (
          nx36160), .B0 (camera_module_cache_ram_159__5), .B1 (nx36200)) ;
    dffr camera_module_cache_reg_ram_143__5 (.Q (camera_module_cache_ram_143__5)
         , .QB (\$dummy [1814]), .D (nx14183), .CLK (clk), .R (rst)) ;
    mux21_ni ix14184 (.Y (nx14183), .A0 (nx35514), .A1 (
             camera_module_cache_ram_143__5), .S0 (nx36760)) ;
    dffr camera_module_cache_reg_ram_159__5 (.Q (camera_module_cache_ram_159__5)
         , .QB (\$dummy [1815]), .D (nx14173), .CLK (clk), .R (rst)) ;
    mux21_ni ix14174 (.Y (nx14173), .A0 (nx35514), .A1 (
             camera_module_cache_ram_159__5), .S0 (nx36764)) ;
    aoi22 ix32217 (.Y (nx32216), .A0 (camera_module_cache_ram_191__5), .A1 (
          nx36240), .B0 (camera_module_cache_ram_175__5), .B1 (nx36280)) ;
    dffr camera_module_cache_reg_ram_191__5 (.Q (camera_module_cache_ram_191__5)
         , .QB (\$dummy [1816]), .D (nx14153), .CLK (clk), .R (rst)) ;
    mux21_ni ix14154 (.Y (nx14153), .A0 (nx35514), .A1 (
             camera_module_cache_ram_191__5), .S0 (nx36768)) ;
    dffr camera_module_cache_reg_ram_175__5 (.Q (camera_module_cache_ram_175__5)
         , .QB (\$dummy [1817]), .D (nx14163), .CLK (clk), .R (rst)) ;
    mux21_ni ix14164 (.Y (nx14163), .A0 (nx35514), .A1 (
             camera_module_cache_ram_175__5), .S0 (nx36772)) ;
    aoi22 ix32225 (.Y (nx32224), .A0 (camera_module_cache_ram_207__5), .A1 (
          nx36320), .B0 (camera_module_cache_ram_223__5), .B1 (nx36360)) ;
    dffr camera_module_cache_reg_ram_207__5 (.Q (camera_module_cache_ram_207__5)
         , .QB (\$dummy [1818]), .D (nx14143), .CLK (clk), .R (rst)) ;
    mux21_ni ix14144 (.Y (nx14143), .A0 (nx35516), .A1 (
             camera_module_cache_ram_207__5), .S0 (nx36776)) ;
    dffr camera_module_cache_reg_ram_223__5 (.Q (camera_module_cache_ram_223__5)
         , .QB (\$dummy [1819]), .D (nx14133), .CLK (clk), .R (rst)) ;
    mux21_ni ix14134 (.Y (nx14133), .A0 (nx35516), .A1 (
             camera_module_cache_ram_223__5), .S0 (nx36780)) ;
    aoi22 ix32233 (.Y (nx32232), .A0 (camera_module_cache_ram_239__5), .A1 (
          nx36400), .B0 (camera_module_cache_ram_255__5), .B1 (nx36440)) ;
    dffr camera_module_cache_reg_ram_239__5 (.Q (camera_module_cache_ram_239__5)
         , .QB (\$dummy [1820]), .D (nx14123), .CLK (clk), .R (rst)) ;
    mux21_ni ix14124 (.Y (nx14123), .A0 (nx35516), .A1 (
             camera_module_cache_ram_239__5), .S0 (nx36784)) ;
    dffr camera_module_cache_reg_ram_255__5 (.Q (camera_module_cache_ram_255__5)
         , .QB (\$dummy [1821]), .D (nx14113), .CLK (clk), .R (rst)) ;
    mux21_ni ix14114 (.Y (nx14113), .A0 (nx35516), .A1 (
             camera_module_cache_ram_255__5), .S0 (nx36788)) ;
    dff camera_module_algo_module_pixel_reg_reg_q_7 (.Q (
        camera_module_algo_module_pixel_value_7), .QB (nx33382), .D (nx21813), .CLK (
        clk)) ;
    mux21_ni ix21814 (.Y (nx21813), .A0 (nx25382), .A1 (
             camera_module_algo_module_pixel_value_7), .S0 (nx22665)) ;
    mux21_ni ix32249 (.Y (nx32248), .A0 (nx32250), .A1 (nx35678), .S0 (nx36794)
             ) ;
    nor04 ix32251 (.Y (nx32250), .A0 (nx25362), .A1 (nx24708), .A2 (nx24052), .A3 (
          nx23398)) ;
    nand04 ix25363 (.Y (nx25362), .A0 (nx32253), .A1 (nx32359), .A2 (nx32427), .A3 (
           nx32495)) ;
    oai21 ix32254 (.Y (nx32253), .A0 (nx25352), .A1 (nx25274), .B0 (nx37232)) ;
    nand04 ix25353 (.Y (nx25352), .A0 (nx32256), .A1 (nx32302), .A2 (nx32310), .A3 (
           nx32318)) ;
    aoi22 ix32257 (.Y (nx32256), .A0 (camera_module_cache_ram_0__7), .A1 (
          nx35840), .B0 (camera_module_cache_ram_16__7), .B1 (nx35880)) ;
    dffr camera_module_cache_reg_ram_0__7 (.Q (camera_module_cache_ram_0__7), .QB (
         \$dummy [1822]), .D (nx21803), .CLK (clk), .R (rst)) ;
    mux21_ni ix21804 (.Y (nx21803), .A0 (camera_module_cache_ram_0__7), .A1 (
             nx35596), .S0 (nx35136)) ;
    oai221 ix22745 (.Y (nx22744), .A0 (nx34076), .A1 (nx32261), .B0 (nx32277), .B1 (
           nx35714), .C0 (nx32280)) ;
    tri01 nvm_module_tri_dataout_127 (.Y (nvm_data_127), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_119 (.Y (nvm_data_119), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_111 (.Y (nvm_data_111), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_103 (.Y (nvm_data_103), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_95 (.Y (nvm_data_95), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_87 (.Y (nvm_data_87), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_79 (.Y (nvm_data_79), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_71 (.Y (nvm_data_71), .A (nx22549), .E (
          nvm_module_GND0)) ;
    inv01 ix32278 (.Y (nx32277), .A (nvm_data_7)) ;
    tri01 nvm_module_tri_dataout_7 (.Y (nvm_data_7), .A (nx22549), .E (
          nvm_module_GND0)) ;
    nand02 ix32281 (.Y (nx32280), .A0 (nx34076), .A1 (nx22678)) ;
    tri01 nvm_module_tri_dataout_63 (.Y (nvm_data_63), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_55 (.Y (nvm_data_55), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_47 (.Y (nvm_data_47), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_39 (.Y (nvm_data_39), .A (nx22549), .E (
          nvm_module_GND0)) ;
    oai22 ix22647 (.Y (nx22646), .A0 (nx34110), .A1 (nx32291), .B0 (nx34096), .B1 (
          nx32295)) ;
    tri01 nvm_module_tri_dataout_31 (.Y (nvm_data_31), .A (nx22549), .E (
          nvm_module_GND0)) ;
    tri01 nvm_module_tri_dataout_23 (.Y (nvm_data_23), .A (nx22549), .E (
          nvm_module_GND0)) ;
    nand02 ix32296 (.Y (nx32295), .A0 (nvm_data_15), .A1 (nx34110)) ;
    tri01 nvm_module_tri_dataout_15 (.Y (nvm_data_15), .A (nx22549), .E (
          nvm_module_GND0)) ;
    dffr camera_module_cache_reg_ram_16__7 (.Q (camera_module_cache_ram_16__7), 
         .QB (\$dummy [1823]), .D (nx21793), .CLK (clk), .R (rst)) ;
    mux21_ni ix21794 (.Y (nx21793), .A0 (camera_module_cache_ram_16__7), .A1 (
             nx35596), .S0 (nx35132)) ;
    aoi22 ix32303 (.Y (nx32302), .A0 (camera_module_cache_ram_32__7), .A1 (
          nx35920), .B0 (camera_module_cache_ram_48__7), .B1 (nx35960)) ;
    dffr camera_module_cache_reg_ram_32__7 (.Q (camera_module_cache_ram_32__7), 
         .QB (\$dummy [1824]), .D (nx21783), .CLK (clk), .R (rst)) ;
    mux21_ni ix21784 (.Y (nx21783), .A0 (camera_module_cache_ram_32__7), .A1 (
             nx35596), .S0 (nx35128)) ;
    dffr camera_module_cache_reg_ram_48__7 (.Q (camera_module_cache_ram_48__7), 
         .QB (\$dummy [1825]), .D (nx21773), .CLK (clk), .R (rst)) ;
    mux21_ni ix21774 (.Y (nx21773), .A0 (camera_module_cache_ram_48__7), .A1 (
             nx35596), .S0 (nx35124)) ;
    aoi22 ix32311 (.Y (nx32310), .A0 (camera_module_cache_ram_64__7), .A1 (
          nx36000), .B0 (camera_module_cache_ram_80__7), .B1 (nx36040)) ;
    dffr camera_module_cache_reg_ram_64__7 (.Q (camera_module_cache_ram_64__7), 
         .QB (\$dummy [1826]), .D (nx21763), .CLK (clk), .R (rst)) ;
    mux21_ni ix21764 (.Y (nx21763), .A0 (camera_module_cache_ram_64__7), .A1 (
             nx35596), .S0 (nx35120)) ;
    dffr camera_module_cache_reg_ram_80__7 (.Q (camera_module_cache_ram_80__7), 
         .QB (\$dummy [1827]), .D (nx21753), .CLK (clk), .R (rst)) ;
    mux21_ni ix21754 (.Y (nx21753), .A0 (camera_module_cache_ram_80__7), .A1 (
             nx35596), .S0 (nx35116)) ;
    aoi22 ix32319 (.Y (nx32318), .A0 (camera_module_cache_ram_112__7), .A1 (
          nx36080), .B0 (camera_module_cache_ram_96__7), .B1 (nx36120)) ;
    dffr camera_module_cache_reg_ram_112__7 (.Q (camera_module_cache_ram_112__7)
         , .QB (\$dummy [1828]), .D (nx21733), .CLK (clk), .R (rst)) ;
    mux21_ni ix21734 (.Y (nx21733), .A0 (camera_module_cache_ram_112__7), .A1 (
             nx35596), .S0 (nx35108)) ;
    dffr camera_module_cache_reg_ram_96__7 (.Q (camera_module_cache_ram_96__7), 
         .QB (\$dummy [1829]), .D (nx21743), .CLK (clk), .R (rst)) ;
    mux21_ni ix21744 (.Y (nx21743), .A0 (camera_module_cache_ram_96__7), .A1 (
             nx35598), .S0 (nx35112)) ;
    nand04 ix25275 (.Y (nx25274), .A0 (nx32327), .A1 (nx32335), .A2 (nx32343), .A3 (
           nx32351)) ;
    aoi22 ix32328 (.Y (nx32327), .A0 (camera_module_cache_ram_128__7), .A1 (
          nx36160), .B0 (camera_module_cache_ram_144__7), .B1 (nx36200)) ;
    dffr camera_module_cache_reg_ram_128__7 (.Q (camera_module_cache_ram_128__7)
         , .QB (\$dummy [1830]), .D (nx21723), .CLK (clk), .R (rst)) ;
    mux21_ni ix21724 (.Y (nx21723), .A0 (camera_module_cache_ram_128__7), .A1 (
             nx35598), .S0 (nx35104)) ;
    dffr camera_module_cache_reg_ram_144__7 (.Q (camera_module_cache_ram_144__7)
         , .QB (\$dummy [1831]), .D (nx21713), .CLK (clk), .R (rst)) ;
    mux21_ni ix21714 (.Y (nx21713), .A0 (camera_module_cache_ram_144__7), .A1 (
             nx35598), .S0 (nx35100)) ;
    aoi22 ix32336 (.Y (nx32335), .A0 (camera_module_cache_ram_176__7), .A1 (
          nx36240), .B0 (camera_module_cache_ram_160__7), .B1 (nx36280)) ;
    dffr camera_module_cache_reg_ram_176__7 (.Q (camera_module_cache_ram_176__7)
         , .QB (\$dummy [1832]), .D (nx21693), .CLK (clk), .R (rst)) ;
    mux21_ni ix21694 (.Y (nx21693), .A0 (camera_module_cache_ram_176__7), .A1 (
             nx35598), .S0 (nx35092)) ;
    dffr camera_module_cache_reg_ram_160__7 (.Q (camera_module_cache_ram_160__7)
         , .QB (\$dummy [1833]), .D (nx21703), .CLK (clk), .R (rst)) ;
    mux21_ni ix21704 (.Y (nx21703), .A0 (camera_module_cache_ram_160__7), .A1 (
             nx35598), .S0 (nx35096)) ;
    aoi22 ix32344 (.Y (nx32343), .A0 (camera_module_cache_ram_192__7), .A1 (
          nx36320), .B0 (camera_module_cache_ram_208__7), .B1 (nx36360)) ;
    dffr camera_module_cache_reg_ram_192__7 (.Q (camera_module_cache_ram_192__7)
         , .QB (\$dummy [1834]), .D (nx21683), .CLK (clk), .R (rst)) ;
    mux21_ni ix21684 (.Y (nx21683), .A0 (camera_module_cache_ram_192__7), .A1 (
             nx35598), .S0 (nx35088)) ;
    dffr camera_module_cache_reg_ram_208__7 (.Q (camera_module_cache_ram_208__7)
         , .QB (\$dummy [1835]), .D (nx21673), .CLK (clk), .R (rst)) ;
    mux21_ni ix21674 (.Y (nx21673), .A0 (camera_module_cache_ram_208__7), .A1 (
             nx35598), .S0 (nx35084)) ;
    aoi22 ix32352 (.Y (nx32351), .A0 (camera_module_cache_ram_224__7), .A1 (
          nx36400), .B0 (camera_module_cache_ram_240__7), .B1 (nx36440)) ;
    dffr camera_module_cache_reg_ram_224__7 (.Q (camera_module_cache_ram_224__7)
         , .QB (\$dummy [1836]), .D (nx21663), .CLK (clk), .R (rst)) ;
    mux21_ni ix21664 (.Y (nx21663), .A0 (camera_module_cache_ram_224__7), .A1 (
             nx35600), .S0 (nx35080)) ;
    dffr camera_module_cache_reg_ram_240__7 (.Q (camera_module_cache_ram_240__7)
         , .QB (\$dummy [1837]), .D (nx21653), .CLK (clk), .R (rst)) ;
    mux21_ni ix21654 (.Y (nx21653), .A0 (camera_module_cache_ram_240__7), .A1 (
             nx35600), .S0 (nx35076)) ;
    oai21 ix32360 (.Y (nx32359), .A0 (nx25190), .A1 (nx25112), .B0 (nx37236)) ;
    nand04 ix25191 (.Y (nx25190), .A0 (nx32362), .A1 (nx32370), .A2 (nx32378), .A3 (
           nx32386)) ;
    aoi22 ix32363 (.Y (nx32362), .A0 (camera_module_cache_ram_1__7), .A1 (
          nx35840), .B0 (camera_module_cache_ram_17__7), .B1 (nx35880)) ;
    dffr camera_module_cache_reg_ram_1__7 (.Q (camera_module_cache_ram_1__7), .QB (
         \$dummy [1838]), .D (nx21643), .CLK (clk), .R (rst)) ;
    mux21_ni ix21644 (.Y (nx21643), .A0 (camera_module_cache_ram_1__7), .A1 (
             nx35600), .S0 (nx35066)) ;
    dffr camera_module_cache_reg_ram_17__7 (.Q (camera_module_cache_ram_17__7), 
         .QB (\$dummy [1839]), .D (nx21633), .CLK (clk), .R (rst)) ;
    mux21_ni ix21634 (.Y (nx21633), .A0 (camera_module_cache_ram_17__7), .A1 (
             nx35600), .S0 (nx35062)) ;
    aoi22 ix32371 (.Y (nx32370), .A0 (camera_module_cache_ram_33__7), .A1 (
          nx35920), .B0 (camera_module_cache_ram_49__7), .B1 (nx35960)) ;
    dffr camera_module_cache_reg_ram_33__7 (.Q (camera_module_cache_ram_33__7), 
         .QB (\$dummy [1840]), .D (nx21623), .CLK (clk), .R (rst)) ;
    mux21_ni ix21624 (.Y (nx21623), .A0 (camera_module_cache_ram_33__7), .A1 (
             nx35600), .S0 (nx35058)) ;
    dffr camera_module_cache_reg_ram_49__7 (.Q (camera_module_cache_ram_49__7), 
         .QB (\$dummy [1841]), .D (nx21613), .CLK (clk), .R (rst)) ;
    mux21_ni ix21614 (.Y (nx21613), .A0 (camera_module_cache_ram_49__7), .A1 (
             nx35600), .S0 (nx35054)) ;
    aoi22 ix32379 (.Y (nx32378), .A0 (camera_module_cache_ram_65__7), .A1 (
          nx36000), .B0 (camera_module_cache_ram_81__7), .B1 (nx36040)) ;
    dffr camera_module_cache_reg_ram_65__7 (.Q (camera_module_cache_ram_65__7), 
         .QB (\$dummy [1842]), .D (nx21603), .CLK (clk), .R (rst)) ;
    mux21_ni ix21604 (.Y (nx21603), .A0 (camera_module_cache_ram_65__7), .A1 (
             nx35600), .S0 (nx35050)) ;
    dffr camera_module_cache_reg_ram_81__7 (.Q (camera_module_cache_ram_81__7), 
         .QB (\$dummy [1843]), .D (nx21593), .CLK (clk), .R (rst)) ;
    mux21_ni ix21594 (.Y (nx21593), .A0 (camera_module_cache_ram_81__7), .A1 (
             nx35602), .S0 (nx35046)) ;
    aoi22 ix32387 (.Y (nx32386), .A0 (camera_module_cache_ram_113__7), .A1 (
          nx36080), .B0 (camera_module_cache_ram_97__7), .B1 (nx36120)) ;
    dffr camera_module_cache_reg_ram_113__7 (.Q (camera_module_cache_ram_113__7)
         , .QB (\$dummy [1844]), .D (nx21573), .CLK (clk), .R (rst)) ;
    mux21_ni ix21574 (.Y (nx21573), .A0 (camera_module_cache_ram_113__7), .A1 (
             nx35602), .S0 (nx35038)) ;
    dffr camera_module_cache_reg_ram_97__7 (.Q (camera_module_cache_ram_97__7), 
         .QB (\$dummy [1845]), .D (nx21583), .CLK (clk), .R (rst)) ;
    mux21_ni ix21584 (.Y (nx21583), .A0 (camera_module_cache_ram_97__7), .A1 (
             nx35602), .S0 (nx35042)) ;
    nand04 ix25113 (.Y (nx25112), .A0 (nx32395), .A1 (nx32403), .A2 (nx32411), .A3 (
           nx32419)) ;
    aoi22 ix32396 (.Y (nx32395), .A0 (camera_module_cache_ram_129__7), .A1 (
          nx36160), .B0 (camera_module_cache_ram_145__7), .B1 (nx36200)) ;
    dffr camera_module_cache_reg_ram_129__7 (.Q (camera_module_cache_ram_129__7)
         , .QB (\$dummy [1846]), .D (nx21563), .CLK (clk), .R (rst)) ;
    mux21_ni ix21564 (.Y (nx21563), .A0 (camera_module_cache_ram_129__7), .A1 (
             nx35602), .S0 (nx35034)) ;
    dffr camera_module_cache_reg_ram_145__7 (.Q (camera_module_cache_ram_145__7)
         , .QB (\$dummy [1847]), .D (nx21553), .CLK (clk), .R (rst)) ;
    mux21_ni ix21554 (.Y (nx21553), .A0 (camera_module_cache_ram_145__7), .A1 (
             nx35602), .S0 (nx35030)) ;
    aoi22 ix32404 (.Y (nx32403), .A0 (camera_module_cache_ram_177__7), .A1 (
          nx36240), .B0 (camera_module_cache_ram_161__7), .B1 (nx36280)) ;
    dffr camera_module_cache_reg_ram_177__7 (.Q (camera_module_cache_ram_177__7)
         , .QB (\$dummy [1848]), .D (nx21533), .CLK (clk), .R (rst)) ;
    mux21_ni ix21534 (.Y (nx21533), .A0 (camera_module_cache_ram_177__7), .A1 (
             nx35602), .S0 (nx35022)) ;
    dffr camera_module_cache_reg_ram_161__7 (.Q (camera_module_cache_ram_161__7)
         , .QB (\$dummy [1849]), .D (nx21543), .CLK (clk), .R (rst)) ;
    mux21_ni ix21544 (.Y (nx21543), .A0 (camera_module_cache_ram_161__7), .A1 (
             nx35602), .S0 (nx35026)) ;
    aoi22 ix32412 (.Y (nx32411), .A0 (camera_module_cache_ram_193__7), .A1 (
          nx36320), .B0 (camera_module_cache_ram_209__7), .B1 (nx36360)) ;
    dffr camera_module_cache_reg_ram_193__7 (.Q (camera_module_cache_ram_193__7)
         , .QB (\$dummy [1850]), .D (nx21523), .CLK (clk), .R (rst)) ;
    mux21_ni ix21524 (.Y (nx21523), .A0 (camera_module_cache_ram_193__7), .A1 (
             nx35604), .S0 (nx35018)) ;
    dffr camera_module_cache_reg_ram_209__7 (.Q (camera_module_cache_ram_209__7)
         , .QB (\$dummy [1851]), .D (nx21513), .CLK (clk), .R (rst)) ;
    mux21_ni ix21514 (.Y (nx21513), .A0 (camera_module_cache_ram_209__7), .A1 (
             nx35604), .S0 (nx35014)) ;
    aoi22 ix32420 (.Y (nx32419), .A0 (camera_module_cache_ram_225__7), .A1 (
          nx36400), .B0 (camera_module_cache_ram_241__7), .B1 (nx36440)) ;
    dffr camera_module_cache_reg_ram_225__7 (.Q (camera_module_cache_ram_225__7)
         , .QB (\$dummy [1852]), .D (nx21503), .CLK (clk), .R (rst)) ;
    mux21_ni ix21504 (.Y (nx21503), .A0 (camera_module_cache_ram_225__7), .A1 (
             nx35604), .S0 (nx35010)) ;
    dffr camera_module_cache_reg_ram_241__7 (.Q (camera_module_cache_ram_241__7)
         , .QB (\$dummy [1853]), .D (nx21493), .CLK (clk), .R (rst)) ;
    mux21_ni ix21494 (.Y (nx21493), .A0 (camera_module_cache_ram_241__7), .A1 (
             nx35604), .S0 (nx35006)) ;
    oai21 ix32428 (.Y (nx32427), .A0 (nx25026), .A1 (nx24948), .B0 (nx37240)) ;
    nand04 ix25027 (.Y (nx25026), .A0 (nx32430), .A1 (nx32438), .A2 (nx32446), .A3 (
           nx32454)) ;
    aoi22 ix32431 (.Y (nx32430), .A0 (camera_module_cache_ram_2__7), .A1 (
          nx35840), .B0 (camera_module_cache_ram_18__7), .B1 (nx35880)) ;
    dffr camera_module_cache_reg_ram_2__7 (.Q (camera_module_cache_ram_2__7), .QB (
         \$dummy [1854]), .D (nx21483), .CLK (clk), .R (rst)) ;
    mux21_ni ix21484 (.Y (nx21483), .A0 (camera_module_cache_ram_2__7), .A1 (
             nx35604), .S0 (nx34996)) ;
    dffr camera_module_cache_reg_ram_18__7 (.Q (camera_module_cache_ram_18__7), 
         .QB (\$dummy [1855]), .D (nx21473), .CLK (clk), .R (rst)) ;
    mux21_ni ix21474 (.Y (nx21473), .A0 (camera_module_cache_ram_18__7), .A1 (
             nx35604), .S0 (nx34992)) ;
    aoi22 ix32439 (.Y (nx32438), .A0 (camera_module_cache_ram_34__7), .A1 (
          nx35920), .B0 (camera_module_cache_ram_50__7), .B1 (nx35960)) ;
    dffr camera_module_cache_reg_ram_34__7 (.Q (camera_module_cache_ram_34__7), 
         .QB (\$dummy [1856]), .D (nx21463), .CLK (clk), .R (rst)) ;
    mux21_ni ix21464 (.Y (nx21463), .A0 (camera_module_cache_ram_34__7), .A1 (
             nx35604), .S0 (nx34988)) ;
    dffr camera_module_cache_reg_ram_50__7 (.Q (camera_module_cache_ram_50__7), 
         .QB (\$dummy [1857]), .D (nx21453), .CLK (clk), .R (rst)) ;
    mux21_ni ix21454 (.Y (nx21453), .A0 (camera_module_cache_ram_50__7), .A1 (
             nx35606), .S0 (nx34984)) ;
    aoi22 ix32447 (.Y (nx32446), .A0 (camera_module_cache_ram_66__7), .A1 (
          nx36000), .B0 (camera_module_cache_ram_82__7), .B1 (nx36040)) ;
    dffr camera_module_cache_reg_ram_66__7 (.Q (camera_module_cache_ram_66__7), 
         .QB (\$dummy [1858]), .D (nx21443), .CLK (clk), .R (rst)) ;
    mux21_ni ix21444 (.Y (nx21443), .A0 (camera_module_cache_ram_66__7), .A1 (
             nx35606), .S0 (nx34980)) ;
    dffr camera_module_cache_reg_ram_82__7 (.Q (camera_module_cache_ram_82__7), 
         .QB (\$dummy [1859]), .D (nx21433), .CLK (clk), .R (rst)) ;
    mux21_ni ix21434 (.Y (nx21433), .A0 (camera_module_cache_ram_82__7), .A1 (
             nx35606), .S0 (nx34976)) ;
    aoi22 ix32455 (.Y (nx32454), .A0 (camera_module_cache_ram_114__7), .A1 (
          nx36080), .B0 (camera_module_cache_ram_98__7), .B1 (nx36120)) ;
    dffr camera_module_cache_reg_ram_114__7 (.Q (camera_module_cache_ram_114__7)
         , .QB (\$dummy [1860]), .D (nx21413), .CLK (clk), .R (rst)) ;
    mux21_ni ix21414 (.Y (nx21413), .A0 (camera_module_cache_ram_114__7), .A1 (
             nx35606), .S0 (nx34968)) ;
    dffr camera_module_cache_reg_ram_98__7 (.Q (camera_module_cache_ram_98__7), 
         .QB (\$dummy [1861]), .D (nx21423), .CLK (clk), .R (rst)) ;
    mux21_ni ix21424 (.Y (nx21423), .A0 (camera_module_cache_ram_98__7), .A1 (
             nx35606), .S0 (nx34972)) ;
    nand04 ix24949 (.Y (nx24948), .A0 (nx32463), .A1 (nx32471), .A2 (nx32479), .A3 (
           nx32487)) ;
    aoi22 ix32464 (.Y (nx32463), .A0 (camera_module_cache_ram_130__7), .A1 (
          nx36160), .B0 (camera_module_cache_ram_146__7), .B1 (nx36200)) ;
    dffr camera_module_cache_reg_ram_130__7 (.Q (camera_module_cache_ram_130__7)
         , .QB (\$dummy [1862]), .D (nx21403), .CLK (clk), .R (rst)) ;
    mux21_ni ix21404 (.Y (nx21403), .A0 (camera_module_cache_ram_130__7), .A1 (
             nx35606), .S0 (nx34964)) ;
    dffr camera_module_cache_reg_ram_146__7 (.Q (camera_module_cache_ram_146__7)
         , .QB (\$dummy [1863]), .D (nx21393), .CLK (clk), .R (rst)) ;
    mux21_ni ix21394 (.Y (nx21393), .A0 (camera_module_cache_ram_146__7), .A1 (
             nx35606), .S0 (nx34960)) ;
    aoi22 ix32472 (.Y (nx32471), .A0 (camera_module_cache_ram_178__7), .A1 (
          nx36240), .B0 (camera_module_cache_ram_162__7), .B1 (nx36280)) ;
    dffr camera_module_cache_reg_ram_178__7 (.Q (camera_module_cache_ram_178__7)
         , .QB (\$dummy [1864]), .D (nx21373), .CLK (clk), .R (rst)) ;
    mux21_ni ix21374 (.Y (nx21373), .A0 (camera_module_cache_ram_178__7), .A1 (
             nx35608), .S0 (nx34952)) ;
    dffr camera_module_cache_reg_ram_162__7 (.Q (camera_module_cache_ram_162__7)
         , .QB (\$dummy [1865]), .D (nx21383), .CLK (clk), .R (rst)) ;
    mux21_ni ix21384 (.Y (nx21383), .A0 (camera_module_cache_ram_162__7), .A1 (
             nx35608), .S0 (nx34956)) ;
    aoi22 ix32480 (.Y (nx32479), .A0 (camera_module_cache_ram_194__7), .A1 (
          nx36320), .B0 (camera_module_cache_ram_210__7), .B1 (nx36360)) ;
    dffr camera_module_cache_reg_ram_194__7 (.Q (camera_module_cache_ram_194__7)
         , .QB (\$dummy [1866]), .D (nx21363), .CLK (clk), .R (rst)) ;
    mux21_ni ix21364 (.Y (nx21363), .A0 (camera_module_cache_ram_194__7), .A1 (
             nx35608), .S0 (nx34948)) ;
    dffr camera_module_cache_reg_ram_210__7 (.Q (camera_module_cache_ram_210__7)
         , .QB (\$dummy [1867]), .D (nx21353), .CLK (clk), .R (rst)) ;
    mux21_ni ix21354 (.Y (nx21353), .A0 (camera_module_cache_ram_210__7), .A1 (
             nx35608), .S0 (nx34944)) ;
    aoi22 ix32488 (.Y (nx32487), .A0 (camera_module_cache_ram_226__7), .A1 (
          nx36400), .B0 (camera_module_cache_ram_242__7), .B1 (nx36440)) ;
    dffr camera_module_cache_reg_ram_226__7 (.Q (camera_module_cache_ram_226__7)
         , .QB (\$dummy [1868]), .D (nx21343), .CLK (clk), .R (rst)) ;
    mux21_ni ix21344 (.Y (nx21343), .A0 (camera_module_cache_ram_226__7), .A1 (
             nx35608), .S0 (nx34940)) ;
    dffr camera_module_cache_reg_ram_242__7 (.Q (camera_module_cache_ram_242__7)
         , .QB (\$dummy [1869]), .D (nx21333), .CLK (clk), .R (rst)) ;
    mux21_ni ix21334 (.Y (nx21333), .A0 (camera_module_cache_ram_242__7), .A1 (
             nx35608), .S0 (nx34936)) ;
    oai21 ix32496 (.Y (nx32495), .A0 (nx24864), .A1 (nx24786), .B0 (nx37244)) ;
    nand04 ix24865 (.Y (nx24864), .A0 (nx32498), .A1 (nx32506), .A2 (nx32514), .A3 (
           nx32522)) ;
    aoi22 ix32499 (.Y (nx32498), .A0 (camera_module_cache_ram_3__7), .A1 (
          nx35842), .B0 (camera_module_cache_ram_19__7), .B1 (nx35882)) ;
    dffr camera_module_cache_reg_ram_3__7 (.Q (camera_module_cache_ram_3__7), .QB (
         \$dummy [1870]), .D (nx21323), .CLK (clk), .R (rst)) ;
    mux21_ni ix21324 (.Y (nx21323), .A0 (camera_module_cache_ram_3__7), .A1 (
             nx35608), .S0 (nx34926)) ;
    dffr camera_module_cache_reg_ram_19__7 (.Q (camera_module_cache_ram_19__7), 
         .QB (\$dummy [1871]), .D (nx21313), .CLK (clk), .R (rst)) ;
    mux21_ni ix21314 (.Y (nx21313), .A0 (camera_module_cache_ram_19__7), .A1 (
             nx35610), .S0 (nx34922)) ;
    aoi22 ix32507 (.Y (nx32506), .A0 (camera_module_cache_ram_35__7), .A1 (
          nx35922), .B0 (camera_module_cache_ram_51__7), .B1 (nx35962)) ;
    dffr camera_module_cache_reg_ram_35__7 (.Q (camera_module_cache_ram_35__7), 
         .QB (\$dummy [1872]), .D (nx21303), .CLK (clk), .R (rst)) ;
    mux21_ni ix21304 (.Y (nx21303), .A0 (camera_module_cache_ram_35__7), .A1 (
             nx35610), .S0 (nx34918)) ;
    dffr camera_module_cache_reg_ram_51__7 (.Q (camera_module_cache_ram_51__7), 
         .QB (\$dummy [1873]), .D (nx21293), .CLK (clk), .R (rst)) ;
    mux21_ni ix21294 (.Y (nx21293), .A0 (camera_module_cache_ram_51__7), .A1 (
             nx35610), .S0 (nx34914)) ;
    aoi22 ix32515 (.Y (nx32514), .A0 (camera_module_cache_ram_67__7), .A1 (
          nx36002), .B0 (camera_module_cache_ram_83__7), .B1 (nx36042)) ;
    dffr camera_module_cache_reg_ram_67__7 (.Q (camera_module_cache_ram_67__7), 
         .QB (\$dummy [1874]), .D (nx21283), .CLK (clk), .R (rst)) ;
    mux21_ni ix21284 (.Y (nx21283), .A0 (camera_module_cache_ram_67__7), .A1 (
             nx35610), .S0 (nx34910)) ;
    dffr camera_module_cache_reg_ram_83__7 (.Q (camera_module_cache_ram_83__7), 
         .QB (\$dummy [1875]), .D (nx21273), .CLK (clk), .R (rst)) ;
    mux21_ni ix21274 (.Y (nx21273), .A0 (camera_module_cache_ram_83__7), .A1 (
             nx35610), .S0 (nx34906)) ;
    aoi22 ix32523 (.Y (nx32522), .A0 (camera_module_cache_ram_115__7), .A1 (
          nx36082), .B0 (camera_module_cache_ram_99__7), .B1 (nx36122)) ;
    dffr camera_module_cache_reg_ram_115__7 (.Q (camera_module_cache_ram_115__7)
         , .QB (\$dummy [1876]), .D (nx21253), .CLK (clk), .R (rst)) ;
    mux21_ni ix21254 (.Y (nx21253), .A0 (camera_module_cache_ram_115__7), .A1 (
             nx35610), .S0 (nx34898)) ;
    dffr camera_module_cache_reg_ram_99__7 (.Q (camera_module_cache_ram_99__7), 
         .QB (\$dummy [1877]), .D (nx21263), .CLK (clk), .R (rst)) ;
    mux21_ni ix21264 (.Y (nx21263), .A0 (camera_module_cache_ram_99__7), .A1 (
             nx35610), .S0 (nx34902)) ;
    nand04 ix24787 (.Y (nx24786), .A0 (nx32531), .A1 (nx32539), .A2 (nx32547), .A3 (
           nx32555)) ;
    aoi22 ix32532 (.Y (nx32531), .A0 (camera_module_cache_ram_131__7), .A1 (
          nx36162), .B0 (camera_module_cache_ram_147__7), .B1 (nx36202)) ;
    dffr camera_module_cache_reg_ram_131__7 (.Q (camera_module_cache_ram_131__7)
         , .QB (\$dummy [1878]), .D (nx21243), .CLK (clk), .R (rst)) ;
    mux21_ni ix21244 (.Y (nx21243), .A0 (camera_module_cache_ram_131__7), .A1 (
             nx35612), .S0 (nx34894)) ;
    dffr camera_module_cache_reg_ram_147__7 (.Q (camera_module_cache_ram_147__7)
         , .QB (\$dummy [1879]), .D (nx21233), .CLK (clk), .R (rst)) ;
    mux21_ni ix21234 (.Y (nx21233), .A0 (camera_module_cache_ram_147__7), .A1 (
             nx35612), .S0 (nx34890)) ;
    aoi22 ix32540 (.Y (nx32539), .A0 (camera_module_cache_ram_179__7), .A1 (
          nx36242), .B0 (camera_module_cache_ram_163__7), .B1 (nx36282)) ;
    dffr camera_module_cache_reg_ram_179__7 (.Q (camera_module_cache_ram_179__7)
         , .QB (\$dummy [1880]), .D (nx21213), .CLK (clk), .R (rst)) ;
    mux21_ni ix21214 (.Y (nx21213), .A0 (camera_module_cache_ram_179__7), .A1 (
             nx35612), .S0 (nx34882)) ;
    dffr camera_module_cache_reg_ram_163__7 (.Q (camera_module_cache_ram_163__7)
         , .QB (\$dummy [1881]), .D (nx21223), .CLK (clk), .R (rst)) ;
    mux21_ni ix21224 (.Y (nx21223), .A0 (camera_module_cache_ram_163__7), .A1 (
             nx35612), .S0 (nx34886)) ;
    aoi22 ix32548 (.Y (nx32547), .A0 (camera_module_cache_ram_195__7), .A1 (
          nx36322), .B0 (camera_module_cache_ram_211__7), .B1 (nx36362)) ;
    dffr camera_module_cache_reg_ram_195__7 (.Q (camera_module_cache_ram_195__7)
         , .QB (\$dummy [1882]), .D (nx21203), .CLK (clk), .R (rst)) ;
    mux21_ni ix21204 (.Y (nx21203), .A0 (camera_module_cache_ram_195__7), .A1 (
             nx35612), .S0 (nx34878)) ;
    dffr camera_module_cache_reg_ram_211__7 (.Q (camera_module_cache_ram_211__7)
         , .QB (\$dummy [1883]), .D (nx21193), .CLK (clk), .R (rst)) ;
    mux21_ni ix21194 (.Y (nx21193), .A0 (camera_module_cache_ram_211__7), .A1 (
             nx35612), .S0 (nx34874)) ;
    aoi22 ix32556 (.Y (nx32555), .A0 (camera_module_cache_ram_227__7), .A1 (
          nx36402), .B0 (camera_module_cache_ram_243__7), .B1 (nx36442)) ;
    dffr camera_module_cache_reg_ram_227__7 (.Q (camera_module_cache_ram_227__7)
         , .QB (\$dummy [1884]), .D (nx21183), .CLK (clk), .R (rst)) ;
    mux21_ni ix21184 (.Y (nx21183), .A0 (camera_module_cache_ram_227__7), .A1 (
             nx35612), .S0 (nx34870)) ;
    dffr camera_module_cache_reg_ram_243__7 (.Q (camera_module_cache_ram_243__7)
         , .QB (\$dummy [1885]), .D (nx21173), .CLK (clk), .R (rst)) ;
    mux21_ni ix21174 (.Y (nx21173), .A0 (camera_module_cache_ram_243__7), .A1 (
             nx35614), .S0 (nx34866)) ;
    nand04 ix24709 (.Y (nx24708), .A0 (nx32564), .A1 (nx32632), .A2 (nx32700), .A3 (
           nx32768)) ;
    oai21 ix32565 (.Y (nx32564), .A0 (nx24698), .A1 (nx24620), .B0 (nx37248)) ;
    nand04 ix24699 (.Y (nx24698), .A0 (nx32567), .A1 (nx32575), .A2 (nx32583), .A3 (
           nx32591)) ;
    aoi22 ix32568 (.Y (nx32567), .A0 (camera_module_cache_ram_4__7), .A1 (
          nx35842), .B0 (camera_module_cache_ram_20__7), .B1 (nx35882)) ;
    dffr camera_module_cache_reg_ram_4__7 (.Q (camera_module_cache_ram_4__7), .QB (
         \$dummy [1886]), .D (nx21163), .CLK (clk), .R (rst)) ;
    mux21_ni ix21164 (.Y (nx21163), .A0 (camera_module_cache_ram_4__7), .A1 (
             nx35614), .S0 (nx34856)) ;
    dffr camera_module_cache_reg_ram_20__7 (.Q (camera_module_cache_ram_20__7), 
         .QB (\$dummy [1887]), .D (nx21153), .CLK (clk), .R (rst)) ;
    mux21_ni ix21154 (.Y (nx21153), .A0 (camera_module_cache_ram_20__7), .A1 (
             nx35614), .S0 (nx34852)) ;
    aoi22 ix32576 (.Y (nx32575), .A0 (camera_module_cache_ram_36__7), .A1 (
          nx35922), .B0 (camera_module_cache_ram_52__7), .B1 (nx35962)) ;
    dffr camera_module_cache_reg_ram_36__7 (.Q (camera_module_cache_ram_36__7), 
         .QB (\$dummy [1888]), .D (nx21143), .CLK (clk), .R (rst)) ;
    mux21_ni ix21144 (.Y (nx21143), .A0 (camera_module_cache_ram_36__7), .A1 (
             nx35614), .S0 (nx34848)) ;
    dffr camera_module_cache_reg_ram_52__7 (.Q (camera_module_cache_ram_52__7), 
         .QB (\$dummy [1889]), .D (nx21133), .CLK (clk), .R (rst)) ;
    mux21_ni ix21134 (.Y (nx21133), .A0 (camera_module_cache_ram_52__7), .A1 (
             nx35614), .S0 (nx34844)) ;
    aoi22 ix32584 (.Y (nx32583), .A0 (camera_module_cache_ram_68__7), .A1 (
          nx36002), .B0 (camera_module_cache_ram_84__7), .B1 (nx36042)) ;
    dffr camera_module_cache_reg_ram_68__7 (.Q (camera_module_cache_ram_68__7), 
         .QB (\$dummy [1890]), .D (nx21123), .CLK (clk), .R (rst)) ;
    mux21_ni ix21124 (.Y (nx21123), .A0 (camera_module_cache_ram_68__7), .A1 (
             nx35614), .S0 (nx34840)) ;
    dffr camera_module_cache_reg_ram_84__7 (.Q (camera_module_cache_ram_84__7), 
         .QB (\$dummy [1891]), .D (nx21113), .CLK (clk), .R (rst)) ;
    mux21_ni ix21114 (.Y (nx21113), .A0 (camera_module_cache_ram_84__7), .A1 (
             nx35614), .S0 (nx34836)) ;
    aoi22 ix32592 (.Y (nx32591), .A0 (camera_module_cache_ram_116__7), .A1 (
          nx36082), .B0 (camera_module_cache_ram_100__7), .B1 (nx36122)) ;
    dffr camera_module_cache_reg_ram_116__7 (.Q (camera_module_cache_ram_116__7)
         , .QB (\$dummy [1892]), .D (nx21093), .CLK (clk), .R (rst)) ;
    mux21_ni ix21094 (.Y (nx21093), .A0 (camera_module_cache_ram_116__7), .A1 (
             nx35616), .S0 (nx34828)) ;
    dffr camera_module_cache_reg_ram_100__7 (.Q (camera_module_cache_ram_100__7)
         , .QB (\$dummy [1893]), .D (nx21103), .CLK (clk), .R (rst)) ;
    mux21_ni ix21104 (.Y (nx21103), .A0 (camera_module_cache_ram_100__7), .A1 (
             nx35616), .S0 (nx34832)) ;
    nand04 ix24621 (.Y (nx24620), .A0 (nx32600), .A1 (nx32608), .A2 (nx32616), .A3 (
           nx32624)) ;
    aoi22 ix32601 (.Y (nx32600), .A0 (camera_module_cache_ram_132__7), .A1 (
          nx36162), .B0 (camera_module_cache_ram_148__7), .B1 (nx36202)) ;
    dffr camera_module_cache_reg_ram_132__7 (.Q (camera_module_cache_ram_132__7)
         , .QB (\$dummy [1894]), .D (nx21083), .CLK (clk), .R (rst)) ;
    mux21_ni ix21084 (.Y (nx21083), .A0 (camera_module_cache_ram_132__7), .A1 (
             nx35616), .S0 (nx34824)) ;
    dffr camera_module_cache_reg_ram_148__7 (.Q (camera_module_cache_ram_148__7)
         , .QB (\$dummy [1895]), .D (nx21073), .CLK (clk), .R (rst)) ;
    mux21_ni ix21074 (.Y (nx21073), .A0 (camera_module_cache_ram_148__7), .A1 (
             nx35616), .S0 (nx34820)) ;
    aoi22 ix32609 (.Y (nx32608), .A0 (camera_module_cache_ram_180__7), .A1 (
          nx36242), .B0 (camera_module_cache_ram_164__7), .B1 (nx36282)) ;
    dffr camera_module_cache_reg_ram_180__7 (.Q (camera_module_cache_ram_180__7)
         , .QB (\$dummy [1896]), .D (nx21053), .CLK (clk), .R (rst)) ;
    mux21_ni ix21054 (.Y (nx21053), .A0 (camera_module_cache_ram_180__7), .A1 (
             nx35616), .S0 (nx34812)) ;
    dffr camera_module_cache_reg_ram_164__7 (.Q (camera_module_cache_ram_164__7)
         , .QB (\$dummy [1897]), .D (nx21063), .CLK (clk), .R (rst)) ;
    mux21_ni ix21064 (.Y (nx21063), .A0 (camera_module_cache_ram_164__7), .A1 (
             nx35616), .S0 (nx34816)) ;
    aoi22 ix32617 (.Y (nx32616), .A0 (camera_module_cache_ram_196__7), .A1 (
          nx36322), .B0 (camera_module_cache_ram_212__7), .B1 (nx36362)) ;
    dffr camera_module_cache_reg_ram_196__7 (.Q (camera_module_cache_ram_196__7)
         , .QB (\$dummy [1898]), .D (nx21043), .CLK (clk), .R (rst)) ;
    mux21_ni ix21044 (.Y (nx21043), .A0 (camera_module_cache_ram_196__7), .A1 (
             nx35616), .S0 (nx34808)) ;
    dffr camera_module_cache_reg_ram_212__7 (.Q (camera_module_cache_ram_212__7)
         , .QB (\$dummy [1899]), .D (nx21033), .CLK (clk), .R (rst)) ;
    mux21_ni ix21034 (.Y (nx21033), .A0 (camera_module_cache_ram_212__7), .A1 (
             nx35618), .S0 (nx34804)) ;
    aoi22 ix32625 (.Y (nx32624), .A0 (camera_module_cache_ram_228__7), .A1 (
          nx36402), .B0 (camera_module_cache_ram_244__7), .B1 (nx36442)) ;
    dffr camera_module_cache_reg_ram_228__7 (.Q (camera_module_cache_ram_228__7)
         , .QB (\$dummy [1900]), .D (nx21023), .CLK (clk), .R (rst)) ;
    mux21_ni ix21024 (.Y (nx21023), .A0 (camera_module_cache_ram_228__7), .A1 (
             nx35618), .S0 (nx34800)) ;
    dffr camera_module_cache_reg_ram_244__7 (.Q (camera_module_cache_ram_244__7)
         , .QB (\$dummy [1901]), .D (nx21013), .CLK (clk), .R (rst)) ;
    mux21_ni ix21014 (.Y (nx21013), .A0 (camera_module_cache_ram_244__7), .A1 (
             nx35618), .S0 (nx34796)) ;
    oai21 ix32633 (.Y (nx32632), .A0 (nx24536), .A1 (nx24458), .B0 (nx37252)) ;
    nand04 ix24537 (.Y (nx24536), .A0 (nx32635), .A1 (nx32643), .A2 (nx32651), .A3 (
           nx32659)) ;
    aoi22 ix32636 (.Y (nx32635), .A0 (camera_module_cache_ram_5__7), .A1 (
          nx35842), .B0 (camera_module_cache_ram_21__7), .B1 (nx35882)) ;
    dffr camera_module_cache_reg_ram_5__7 (.Q (camera_module_cache_ram_5__7), .QB (
         \$dummy [1902]), .D (nx21003), .CLK (clk), .R (rst)) ;
    mux21_ni ix21004 (.Y (nx21003), .A0 (camera_module_cache_ram_5__7), .A1 (
             nx35618), .S0 (nx34786)) ;
    dffr camera_module_cache_reg_ram_21__7 (.Q (camera_module_cache_ram_21__7), 
         .QB (\$dummy [1903]), .D (nx20993), .CLK (clk), .R (rst)) ;
    mux21_ni ix20994 (.Y (nx20993), .A0 (camera_module_cache_ram_21__7), .A1 (
             nx35618), .S0 (nx34782)) ;
    aoi22 ix32644 (.Y (nx32643), .A0 (camera_module_cache_ram_37__7), .A1 (
          nx35922), .B0 (camera_module_cache_ram_53__7), .B1 (nx35962)) ;
    dffr camera_module_cache_reg_ram_37__7 (.Q (camera_module_cache_ram_37__7), 
         .QB (\$dummy [1904]), .D (nx20983), .CLK (clk), .R (rst)) ;
    mux21_ni ix20984 (.Y (nx20983), .A0 (camera_module_cache_ram_37__7), .A1 (
             nx35618), .S0 (nx34778)) ;
    dffr camera_module_cache_reg_ram_53__7 (.Q (camera_module_cache_ram_53__7), 
         .QB (\$dummy [1905]), .D (nx20973), .CLK (clk), .R (rst)) ;
    mux21_ni ix20974 (.Y (nx20973), .A0 (camera_module_cache_ram_53__7), .A1 (
             nx35618), .S0 (nx34774)) ;
    aoi22 ix32652 (.Y (nx32651), .A0 (camera_module_cache_ram_69__7), .A1 (
          nx36002), .B0 (camera_module_cache_ram_85__7), .B1 (nx36042)) ;
    dffr camera_module_cache_reg_ram_69__7 (.Q (camera_module_cache_ram_69__7), 
         .QB (\$dummy [1906]), .D (nx20963), .CLK (clk), .R (rst)) ;
    mux21_ni ix20964 (.Y (nx20963), .A0 (camera_module_cache_ram_69__7), .A1 (
             nx35620), .S0 (nx34770)) ;
    dffr camera_module_cache_reg_ram_85__7 (.Q (camera_module_cache_ram_85__7), 
         .QB (\$dummy [1907]), .D (nx20953), .CLK (clk), .R (rst)) ;
    mux21_ni ix20954 (.Y (nx20953), .A0 (camera_module_cache_ram_85__7), .A1 (
             nx35620), .S0 (nx34766)) ;
    aoi22 ix32660 (.Y (nx32659), .A0 (camera_module_cache_ram_117__7), .A1 (
          nx36082), .B0 (camera_module_cache_ram_101__7), .B1 (nx36122)) ;
    dffr camera_module_cache_reg_ram_117__7 (.Q (camera_module_cache_ram_117__7)
         , .QB (\$dummy [1908]), .D (nx20933), .CLK (clk), .R (rst)) ;
    mux21_ni ix20934 (.Y (nx20933), .A0 (camera_module_cache_ram_117__7), .A1 (
             nx35620), .S0 (nx34758)) ;
    dffr camera_module_cache_reg_ram_101__7 (.Q (camera_module_cache_ram_101__7)
         , .QB (\$dummy [1909]), .D (nx20943), .CLK (clk), .R (rst)) ;
    mux21_ni ix20944 (.Y (nx20943), .A0 (camera_module_cache_ram_101__7), .A1 (
             nx35620), .S0 (nx34762)) ;
    nand04 ix24459 (.Y (nx24458), .A0 (nx32668), .A1 (nx32676), .A2 (nx32684), .A3 (
           nx32692)) ;
    aoi22 ix32669 (.Y (nx32668), .A0 (camera_module_cache_ram_133__7), .A1 (
          nx36162), .B0 (camera_module_cache_ram_149__7), .B1 (nx36202)) ;
    dffr camera_module_cache_reg_ram_133__7 (.Q (camera_module_cache_ram_133__7)
         , .QB (\$dummy [1910]), .D (nx20923), .CLK (clk), .R (rst)) ;
    mux21_ni ix20924 (.Y (nx20923), .A0 (camera_module_cache_ram_133__7), .A1 (
             nx35620), .S0 (nx34754)) ;
    dffr camera_module_cache_reg_ram_149__7 (.Q (camera_module_cache_ram_149__7)
         , .QB (\$dummy [1911]), .D (nx20913), .CLK (clk), .R (rst)) ;
    mux21_ni ix20914 (.Y (nx20913), .A0 (camera_module_cache_ram_149__7), .A1 (
             nx35620), .S0 (nx34750)) ;
    aoi22 ix32677 (.Y (nx32676), .A0 (camera_module_cache_ram_181__7), .A1 (
          nx36242), .B0 (camera_module_cache_ram_165__7), .B1 (nx36282)) ;
    dffr camera_module_cache_reg_ram_181__7 (.Q (camera_module_cache_ram_181__7)
         , .QB (\$dummy [1912]), .D (nx20893), .CLK (clk), .R (rst)) ;
    mux21_ni ix20894 (.Y (nx20893), .A0 (camera_module_cache_ram_181__7), .A1 (
             nx35620), .S0 (nx34742)) ;
    dffr camera_module_cache_reg_ram_165__7 (.Q (camera_module_cache_ram_165__7)
         , .QB (\$dummy [1913]), .D (nx20903), .CLK (clk), .R (rst)) ;
    mux21_ni ix20904 (.Y (nx20903), .A0 (camera_module_cache_ram_165__7), .A1 (
             nx35622), .S0 (nx34746)) ;
    aoi22 ix32685 (.Y (nx32684), .A0 (camera_module_cache_ram_197__7), .A1 (
          nx36322), .B0 (camera_module_cache_ram_213__7), .B1 (nx36362)) ;
    dffr camera_module_cache_reg_ram_197__7 (.Q (camera_module_cache_ram_197__7)
         , .QB (\$dummy [1914]), .D (nx20883), .CLK (clk), .R (rst)) ;
    mux21_ni ix20884 (.Y (nx20883), .A0 (camera_module_cache_ram_197__7), .A1 (
             nx35622), .S0 (nx34738)) ;
    dffr camera_module_cache_reg_ram_213__7 (.Q (camera_module_cache_ram_213__7)
         , .QB (\$dummy [1915]), .D (nx20873), .CLK (clk), .R (rst)) ;
    mux21_ni ix20874 (.Y (nx20873), .A0 (camera_module_cache_ram_213__7), .A1 (
             nx35622), .S0 (nx34734)) ;
    aoi22 ix32693 (.Y (nx32692), .A0 (camera_module_cache_ram_229__7), .A1 (
          nx36402), .B0 (camera_module_cache_ram_245__7), .B1 (nx36442)) ;
    dffr camera_module_cache_reg_ram_229__7 (.Q (camera_module_cache_ram_229__7)
         , .QB (\$dummy [1916]), .D (nx20863), .CLK (clk), .R (rst)) ;
    mux21_ni ix20864 (.Y (nx20863), .A0 (camera_module_cache_ram_229__7), .A1 (
             nx35622), .S0 (nx34730)) ;
    dffr camera_module_cache_reg_ram_245__7 (.Q (camera_module_cache_ram_245__7)
         , .QB (\$dummy [1917]), .D (nx20853), .CLK (clk), .R (rst)) ;
    mux21_ni ix20854 (.Y (nx20853), .A0 (camera_module_cache_ram_245__7), .A1 (
             nx35622), .S0 (nx34726)) ;
    oai21 ix32701 (.Y (nx32700), .A0 (nx24372), .A1 (nx24294), .B0 (nx37256)) ;
    nand04 ix24373 (.Y (nx24372), .A0 (nx32703), .A1 (nx32711), .A2 (nx32719), .A3 (
           nx32727)) ;
    aoi22 ix32704 (.Y (nx32703), .A0 (camera_module_cache_ram_6__7), .A1 (
          nx35842), .B0 (camera_module_cache_ram_22__7), .B1 (nx35882)) ;
    dffr camera_module_cache_reg_ram_6__7 (.Q (camera_module_cache_ram_6__7), .QB (
         \$dummy [1918]), .D (nx20843), .CLK (clk), .R (rst)) ;
    mux21_ni ix20844 (.Y (nx20843), .A0 (camera_module_cache_ram_6__7), .A1 (
             nx35622), .S0 (nx34716)) ;
    dffr camera_module_cache_reg_ram_22__7 (.Q (camera_module_cache_ram_22__7), 
         .QB (\$dummy [1919]), .D (nx20833), .CLK (clk), .R (rst)) ;
    mux21_ni ix20834 (.Y (nx20833), .A0 (camera_module_cache_ram_22__7), .A1 (
             nx35622), .S0 (nx34712)) ;
    aoi22 ix32712 (.Y (nx32711), .A0 (camera_module_cache_ram_38__7), .A1 (
          nx35922), .B0 (camera_module_cache_ram_54__7), .B1 (nx35962)) ;
    dffr camera_module_cache_reg_ram_38__7 (.Q (camera_module_cache_ram_38__7), 
         .QB (\$dummy [1920]), .D (nx20823), .CLK (clk), .R (rst)) ;
    mux21_ni ix20824 (.Y (nx20823), .A0 (camera_module_cache_ram_38__7), .A1 (
             nx35624), .S0 (nx34708)) ;
    dffr camera_module_cache_reg_ram_54__7 (.Q (camera_module_cache_ram_54__7), 
         .QB (\$dummy [1921]), .D (nx20813), .CLK (clk), .R (rst)) ;
    mux21_ni ix20814 (.Y (nx20813), .A0 (camera_module_cache_ram_54__7), .A1 (
             nx35624), .S0 (nx34704)) ;
    aoi22 ix32720 (.Y (nx32719), .A0 (camera_module_cache_ram_70__7), .A1 (
          nx36002), .B0 (camera_module_cache_ram_86__7), .B1 (nx36042)) ;
    dffr camera_module_cache_reg_ram_70__7 (.Q (camera_module_cache_ram_70__7), 
         .QB (\$dummy [1922]), .D (nx20803), .CLK (clk), .R (rst)) ;
    mux21_ni ix20804 (.Y (nx20803), .A0 (camera_module_cache_ram_70__7), .A1 (
             nx35624), .S0 (nx34700)) ;
    dffr camera_module_cache_reg_ram_86__7 (.Q (camera_module_cache_ram_86__7), 
         .QB (\$dummy [1923]), .D (nx20793), .CLK (clk), .R (rst)) ;
    mux21_ni ix20794 (.Y (nx20793), .A0 (camera_module_cache_ram_86__7), .A1 (
             nx35624), .S0 (nx34696)) ;
    aoi22 ix32728 (.Y (nx32727), .A0 (camera_module_cache_ram_118__7), .A1 (
          nx36082), .B0 (camera_module_cache_ram_102__7), .B1 (nx36122)) ;
    dffr camera_module_cache_reg_ram_118__7 (.Q (camera_module_cache_ram_118__7)
         , .QB (\$dummy [1924]), .D (nx20773), .CLK (clk), .R (rst)) ;
    mux21_ni ix20774 (.Y (nx20773), .A0 (camera_module_cache_ram_118__7), .A1 (
             nx35624), .S0 (nx34688)) ;
    dffr camera_module_cache_reg_ram_102__7 (.Q (camera_module_cache_ram_102__7)
         , .QB (\$dummy [1925]), .D (nx20783), .CLK (clk), .R (rst)) ;
    mux21_ni ix20784 (.Y (nx20783), .A0 (camera_module_cache_ram_102__7), .A1 (
             nx35624), .S0 (nx34692)) ;
    nand04 ix24295 (.Y (nx24294), .A0 (nx32736), .A1 (nx32744), .A2 (nx32752), .A3 (
           nx32760)) ;
    aoi22 ix32737 (.Y (nx32736), .A0 (camera_module_cache_ram_134__7), .A1 (
          nx36162), .B0 (camera_module_cache_ram_150__7), .B1 (nx36202)) ;
    dffr camera_module_cache_reg_ram_134__7 (.Q (camera_module_cache_ram_134__7)
         , .QB (\$dummy [1926]), .D (nx20763), .CLK (clk), .R (rst)) ;
    mux21_ni ix20764 (.Y (nx20763), .A0 (camera_module_cache_ram_134__7), .A1 (
             nx35624), .S0 (nx34684)) ;
    dffr camera_module_cache_reg_ram_150__7 (.Q (camera_module_cache_ram_150__7)
         , .QB (\$dummy [1927]), .D (nx20753), .CLK (clk), .R (rst)) ;
    mux21_ni ix20754 (.Y (nx20753), .A0 (camera_module_cache_ram_150__7), .A1 (
             nx35626), .S0 (nx34680)) ;
    aoi22 ix32745 (.Y (nx32744), .A0 (camera_module_cache_ram_182__7), .A1 (
          nx36242), .B0 (camera_module_cache_ram_166__7), .B1 (nx36282)) ;
    dffr camera_module_cache_reg_ram_182__7 (.Q (camera_module_cache_ram_182__7)
         , .QB (\$dummy [1928]), .D (nx20733), .CLK (clk), .R (rst)) ;
    mux21_ni ix20734 (.Y (nx20733), .A0 (camera_module_cache_ram_182__7), .A1 (
             nx35626), .S0 (nx34672)) ;
    dffr camera_module_cache_reg_ram_166__7 (.Q (camera_module_cache_ram_166__7)
         , .QB (\$dummy [1929]), .D (nx20743), .CLK (clk), .R (rst)) ;
    mux21_ni ix20744 (.Y (nx20743), .A0 (camera_module_cache_ram_166__7), .A1 (
             nx35626), .S0 (nx34676)) ;
    aoi22 ix32753 (.Y (nx32752), .A0 (camera_module_cache_ram_198__7), .A1 (
          nx36322), .B0 (camera_module_cache_ram_214__7), .B1 (nx36362)) ;
    dffr camera_module_cache_reg_ram_198__7 (.Q (camera_module_cache_ram_198__7)
         , .QB (\$dummy [1930]), .D (nx20723), .CLK (clk), .R (rst)) ;
    mux21_ni ix20724 (.Y (nx20723), .A0 (camera_module_cache_ram_198__7), .A1 (
             nx35626), .S0 (nx34668)) ;
    dffr camera_module_cache_reg_ram_214__7 (.Q (camera_module_cache_ram_214__7)
         , .QB (\$dummy [1931]), .D (nx20713), .CLK (clk), .R (rst)) ;
    mux21_ni ix20714 (.Y (nx20713), .A0 (camera_module_cache_ram_214__7), .A1 (
             nx35626), .S0 (nx34664)) ;
    aoi22 ix32761 (.Y (nx32760), .A0 (camera_module_cache_ram_230__7), .A1 (
          nx36402), .B0 (camera_module_cache_ram_246__7), .B1 (nx36442)) ;
    dffr camera_module_cache_reg_ram_230__7 (.Q (camera_module_cache_ram_230__7)
         , .QB (\$dummy [1932]), .D (nx20703), .CLK (clk), .R (rst)) ;
    mux21_ni ix20704 (.Y (nx20703), .A0 (camera_module_cache_ram_230__7), .A1 (
             nx35626), .S0 (nx34660)) ;
    dffr camera_module_cache_reg_ram_246__7 (.Q (camera_module_cache_ram_246__7)
         , .QB (\$dummy [1933]), .D (nx20693), .CLK (clk), .R (rst)) ;
    mux21_ni ix20694 (.Y (nx20693), .A0 (camera_module_cache_ram_246__7), .A1 (
             nx35626), .S0 (nx34656)) ;
    oai21 ix32769 (.Y (nx32768), .A0 (nx24210), .A1 (nx24132), .B0 (nx37260)) ;
    nand04 ix24211 (.Y (nx24210), .A0 (nx32771), .A1 (nx32779), .A2 (nx32787), .A3 (
           nx32795)) ;
    aoi22 ix32772 (.Y (nx32771), .A0 (camera_module_cache_ram_7__7), .A1 (
          nx35842), .B0 (camera_module_cache_ram_23__7), .B1 (nx35882)) ;
    dffr camera_module_cache_reg_ram_7__7 (.Q (camera_module_cache_ram_7__7), .QB (
         \$dummy [1934]), .D (nx20683), .CLK (clk), .R (rst)) ;
    mux21_ni ix20684 (.Y (nx20683), .A0 (camera_module_cache_ram_7__7), .A1 (
             nx35628), .S0 (nx34646)) ;
    dffr camera_module_cache_reg_ram_23__7 (.Q (camera_module_cache_ram_23__7), 
         .QB (\$dummy [1935]), .D (nx20673), .CLK (clk), .R (rst)) ;
    mux21_ni ix20674 (.Y (nx20673), .A0 (camera_module_cache_ram_23__7), .A1 (
             nx35628), .S0 (nx34642)) ;
    aoi22 ix32780 (.Y (nx32779), .A0 (camera_module_cache_ram_39__7), .A1 (
          nx35922), .B0 (camera_module_cache_ram_55__7), .B1 (nx35962)) ;
    dffr camera_module_cache_reg_ram_39__7 (.Q (camera_module_cache_ram_39__7), 
         .QB (\$dummy [1936]), .D (nx20663), .CLK (clk), .R (rst)) ;
    mux21_ni ix20664 (.Y (nx20663), .A0 (camera_module_cache_ram_39__7), .A1 (
             nx35628), .S0 (nx34638)) ;
    dffr camera_module_cache_reg_ram_55__7 (.Q (camera_module_cache_ram_55__7), 
         .QB (\$dummy [1937]), .D (nx20653), .CLK (clk), .R (rst)) ;
    mux21_ni ix20654 (.Y (nx20653), .A0 (camera_module_cache_ram_55__7), .A1 (
             nx35628), .S0 (nx34634)) ;
    aoi22 ix32788 (.Y (nx32787), .A0 (camera_module_cache_ram_71__7), .A1 (
          nx36002), .B0 (camera_module_cache_ram_87__7), .B1 (nx36042)) ;
    dffr camera_module_cache_reg_ram_71__7 (.Q (camera_module_cache_ram_71__7), 
         .QB (\$dummy [1938]), .D (nx20643), .CLK (clk), .R (rst)) ;
    mux21_ni ix20644 (.Y (nx20643), .A0 (camera_module_cache_ram_71__7), .A1 (
             nx35628), .S0 (nx34630)) ;
    dffr camera_module_cache_reg_ram_87__7 (.Q (camera_module_cache_ram_87__7), 
         .QB (\$dummy [1939]), .D (nx20633), .CLK (clk), .R (rst)) ;
    mux21_ni ix20634 (.Y (nx20633), .A0 (camera_module_cache_ram_87__7), .A1 (
             nx35628), .S0 (nx34626)) ;
    aoi22 ix32796 (.Y (nx32795), .A0 (camera_module_cache_ram_119__7), .A1 (
          nx36082), .B0 (camera_module_cache_ram_103__7), .B1 (nx36122)) ;
    dffr camera_module_cache_reg_ram_119__7 (.Q (camera_module_cache_ram_119__7)
         , .QB (\$dummy [1940]), .D (nx20613), .CLK (clk), .R (rst)) ;
    mux21_ni ix20614 (.Y (nx20613), .A0 (camera_module_cache_ram_119__7), .A1 (
             nx35628), .S0 (nx34618)) ;
    dffr camera_module_cache_reg_ram_103__7 (.Q (camera_module_cache_ram_103__7)
         , .QB (\$dummy [1941]), .D (nx20623), .CLK (clk), .R (rst)) ;
    mux21_ni ix20624 (.Y (nx20623), .A0 (camera_module_cache_ram_103__7), .A1 (
             nx35630), .S0 (nx34622)) ;
    nand04 ix24133 (.Y (nx24132), .A0 (nx32804), .A1 (nx32812), .A2 (nx32820), .A3 (
           nx32828)) ;
    aoi22 ix32805 (.Y (nx32804), .A0 (camera_module_cache_ram_135__7), .A1 (
          nx36162), .B0 (camera_module_cache_ram_151__7), .B1 (nx36202)) ;
    dffr camera_module_cache_reg_ram_135__7 (.Q (camera_module_cache_ram_135__7)
         , .QB (\$dummy [1942]), .D (nx20603), .CLK (clk), .R (rst)) ;
    mux21_ni ix20604 (.Y (nx20603), .A0 (camera_module_cache_ram_135__7), .A1 (
             nx35630), .S0 (nx34614)) ;
    dffr camera_module_cache_reg_ram_151__7 (.Q (camera_module_cache_ram_151__7)
         , .QB (\$dummy [1943]), .D (nx20593), .CLK (clk), .R (rst)) ;
    mux21_ni ix20594 (.Y (nx20593), .A0 (camera_module_cache_ram_151__7), .A1 (
             nx35630), .S0 (nx34610)) ;
    aoi22 ix32813 (.Y (nx32812), .A0 (camera_module_cache_ram_183__7), .A1 (
          nx36242), .B0 (camera_module_cache_ram_167__7), .B1 (nx36282)) ;
    dffr camera_module_cache_reg_ram_183__7 (.Q (camera_module_cache_ram_183__7)
         , .QB (\$dummy [1944]), .D (nx20573), .CLK (clk), .R (rst)) ;
    mux21_ni ix20574 (.Y (nx20573), .A0 (camera_module_cache_ram_183__7), .A1 (
             nx35630), .S0 (nx34602)) ;
    dffr camera_module_cache_reg_ram_167__7 (.Q (camera_module_cache_ram_167__7)
         , .QB (\$dummy [1945]), .D (nx20583), .CLK (clk), .R (rst)) ;
    mux21_ni ix20584 (.Y (nx20583), .A0 (camera_module_cache_ram_167__7), .A1 (
             nx35630), .S0 (nx34606)) ;
    aoi22 ix32821 (.Y (nx32820), .A0 (camera_module_cache_ram_199__7), .A1 (
          nx36322), .B0 (camera_module_cache_ram_215__7), .B1 (nx36362)) ;
    dffr camera_module_cache_reg_ram_199__7 (.Q (camera_module_cache_ram_199__7)
         , .QB (\$dummy [1946]), .D (nx20563), .CLK (clk), .R (rst)) ;
    mux21_ni ix20564 (.Y (nx20563), .A0 (camera_module_cache_ram_199__7), .A1 (
             nx35630), .S0 (nx34598)) ;
    dffr camera_module_cache_reg_ram_215__7 (.Q (camera_module_cache_ram_215__7)
         , .QB (\$dummy [1947]), .D (nx20553), .CLK (clk), .R (rst)) ;
    mux21_ni ix20554 (.Y (nx20553), .A0 (camera_module_cache_ram_215__7), .A1 (
             nx35630), .S0 (nx34594)) ;
    aoi22 ix32829 (.Y (nx32828), .A0 (camera_module_cache_ram_231__7), .A1 (
          nx36402), .B0 (camera_module_cache_ram_247__7), .B1 (nx36442)) ;
    dffr camera_module_cache_reg_ram_231__7 (.Q (camera_module_cache_ram_231__7)
         , .QB (\$dummy [1948]), .D (nx20543), .CLK (clk), .R (rst)) ;
    mux21_ni ix20544 (.Y (nx20543), .A0 (camera_module_cache_ram_231__7), .A1 (
             nx35632), .S0 (nx34590)) ;
    dffr camera_module_cache_reg_ram_247__7 (.Q (camera_module_cache_ram_247__7)
         , .QB (\$dummy [1949]), .D (nx20533), .CLK (clk), .R (rst)) ;
    mux21_ni ix20534 (.Y (nx20533), .A0 (camera_module_cache_ram_247__7), .A1 (
             nx35632), .S0 (nx34586)) ;
    nand04 ix24053 (.Y (nx24052), .A0 (nx32837), .A1 (nx32905), .A2 (nx32973), .A3 (
           nx33041)) ;
    oai21 ix32838 (.Y (nx32837), .A0 (nx24042), .A1 (nx23964), .B0 (nx37264)) ;
    nand04 ix24043 (.Y (nx24042), .A0 (nx32840), .A1 (nx32848), .A2 (nx32856), .A3 (
           nx32864)) ;
    aoi22 ix32841 (.Y (nx32840), .A0 (camera_module_cache_ram_8__7), .A1 (
          nx35842), .B0 (camera_module_cache_ram_24__7), .B1 (nx35882)) ;
    dffr camera_module_cache_reg_ram_8__7 (.Q (camera_module_cache_ram_8__7), .QB (
         \$dummy [1950]), .D (nx20523), .CLK (clk), .R (rst)) ;
    mux21_ni ix20524 (.Y (nx20523), .A0 (camera_module_cache_ram_8__7), .A1 (
             nx35632), .S0 (nx34576)) ;
    dffr camera_module_cache_reg_ram_24__7 (.Q (camera_module_cache_ram_24__7), 
         .QB (\$dummy [1951]), .D (nx20513), .CLK (clk), .R (rst)) ;
    mux21_ni ix20514 (.Y (nx20513), .A0 (camera_module_cache_ram_24__7), .A1 (
             nx35632), .S0 (nx34572)) ;
    aoi22 ix32849 (.Y (nx32848), .A0 (camera_module_cache_ram_40__7), .A1 (
          nx35922), .B0 (camera_module_cache_ram_56__7), .B1 (nx35962)) ;
    dffr camera_module_cache_reg_ram_40__7 (.Q (camera_module_cache_ram_40__7), 
         .QB (\$dummy [1952]), .D (nx20503), .CLK (clk), .R (rst)) ;
    mux21_ni ix20504 (.Y (nx20503), .A0 (camera_module_cache_ram_40__7), .A1 (
             nx35632), .S0 (nx34568)) ;
    dffr camera_module_cache_reg_ram_56__7 (.Q (camera_module_cache_ram_56__7), 
         .QB (\$dummy [1953]), .D (nx20493), .CLK (clk), .R (rst)) ;
    mux21_ni ix20494 (.Y (nx20493), .A0 (camera_module_cache_ram_56__7), .A1 (
             nx35632), .S0 (nx34564)) ;
    aoi22 ix32857 (.Y (nx32856), .A0 (camera_module_cache_ram_72__7), .A1 (
          nx36002), .B0 (camera_module_cache_ram_88__7), .B1 (nx36042)) ;
    dffr camera_module_cache_reg_ram_72__7 (.Q (camera_module_cache_ram_72__7), 
         .QB (\$dummy [1954]), .D (nx20483), .CLK (clk), .R (rst)) ;
    mux21_ni ix20484 (.Y (nx20483), .A0 (camera_module_cache_ram_72__7), .A1 (
             nx35632), .S0 (nx34560)) ;
    dffr camera_module_cache_reg_ram_88__7 (.Q (camera_module_cache_ram_88__7), 
         .QB (\$dummy [1955]), .D (nx20473), .CLK (clk), .R (rst)) ;
    mux21_ni ix20474 (.Y (nx20473), .A0 (camera_module_cache_ram_88__7), .A1 (
             nx35634), .S0 (nx34556)) ;
    aoi22 ix32865 (.Y (nx32864), .A0 (camera_module_cache_ram_120__7), .A1 (
          nx36082), .B0 (camera_module_cache_ram_104__7), .B1 (nx36122)) ;
    dffr camera_module_cache_reg_ram_120__7 (.Q (camera_module_cache_ram_120__7)
         , .QB (\$dummy [1956]), .D (nx20453), .CLK (clk), .R (rst)) ;
    mux21_ni ix20454 (.Y (nx20453), .A0 (camera_module_cache_ram_120__7), .A1 (
             nx35634), .S0 (nx34548)) ;
    dffr camera_module_cache_reg_ram_104__7 (.Q (camera_module_cache_ram_104__7)
         , .QB (\$dummy [1957]), .D (nx20463), .CLK (clk), .R (rst)) ;
    mux21_ni ix20464 (.Y (nx20463), .A0 (camera_module_cache_ram_104__7), .A1 (
             nx35634), .S0 (nx34552)) ;
    nand04 ix23965 (.Y (nx23964), .A0 (nx32873), .A1 (nx32881), .A2 (nx32889), .A3 (
           nx32897)) ;
    aoi22 ix32874 (.Y (nx32873), .A0 (camera_module_cache_ram_136__7), .A1 (
          nx36162), .B0 (camera_module_cache_ram_152__7), .B1 (nx36202)) ;
    dffr camera_module_cache_reg_ram_136__7 (.Q (camera_module_cache_ram_136__7)
         , .QB (\$dummy [1958]), .D (nx20443), .CLK (clk), .R (rst)) ;
    mux21_ni ix20444 (.Y (nx20443), .A0 (camera_module_cache_ram_136__7), .A1 (
             nx35634), .S0 (nx34544)) ;
    dffr camera_module_cache_reg_ram_152__7 (.Q (camera_module_cache_ram_152__7)
         , .QB (\$dummy [1959]), .D (nx20433), .CLK (clk), .R (rst)) ;
    mux21_ni ix20434 (.Y (nx20433), .A0 (camera_module_cache_ram_152__7), .A1 (
             nx35634), .S0 (nx34540)) ;
    aoi22 ix32882 (.Y (nx32881), .A0 (camera_module_cache_ram_184__7), .A1 (
          nx36242), .B0 (camera_module_cache_ram_168__7), .B1 (nx36282)) ;
    dffr camera_module_cache_reg_ram_184__7 (.Q (camera_module_cache_ram_184__7)
         , .QB (\$dummy [1960]), .D (nx20413), .CLK (clk), .R (rst)) ;
    mux21_ni ix20414 (.Y (nx20413), .A0 (camera_module_cache_ram_184__7), .A1 (
             nx35634), .S0 (nx34532)) ;
    dffr camera_module_cache_reg_ram_168__7 (.Q (camera_module_cache_ram_168__7)
         , .QB (\$dummy [1961]), .D (nx20423), .CLK (clk), .R (rst)) ;
    mux21_ni ix20424 (.Y (nx20423), .A0 (camera_module_cache_ram_168__7), .A1 (
             nx35634), .S0 (nx34536)) ;
    aoi22 ix32890 (.Y (nx32889), .A0 (camera_module_cache_ram_200__7), .A1 (
          nx36322), .B0 (camera_module_cache_ram_216__7), .B1 (nx36362)) ;
    dffr camera_module_cache_reg_ram_200__7 (.Q (camera_module_cache_ram_200__7)
         , .QB (\$dummy [1962]), .D (nx20403), .CLK (clk), .R (rst)) ;
    mux21_ni ix20404 (.Y (nx20403), .A0 (camera_module_cache_ram_200__7), .A1 (
             nx35636), .S0 (nx34528)) ;
    dffr camera_module_cache_reg_ram_216__7 (.Q (camera_module_cache_ram_216__7)
         , .QB (\$dummy [1963]), .D (nx20393), .CLK (clk), .R (rst)) ;
    mux21_ni ix20394 (.Y (nx20393), .A0 (camera_module_cache_ram_216__7), .A1 (
             nx35636), .S0 (nx34524)) ;
    aoi22 ix32898 (.Y (nx32897), .A0 (camera_module_cache_ram_232__7), .A1 (
          nx36402), .B0 (camera_module_cache_ram_248__7), .B1 (nx36442)) ;
    dffr camera_module_cache_reg_ram_232__7 (.Q (camera_module_cache_ram_232__7)
         , .QB (\$dummy [1964]), .D (nx20383), .CLK (clk), .R (rst)) ;
    mux21_ni ix20384 (.Y (nx20383), .A0 (camera_module_cache_ram_232__7), .A1 (
             nx35636), .S0 (nx34520)) ;
    dffr camera_module_cache_reg_ram_248__7 (.Q (camera_module_cache_ram_248__7)
         , .QB (\$dummy [1965]), .D (nx20373), .CLK (clk), .R (rst)) ;
    mux21_ni ix20374 (.Y (nx20373), .A0 (camera_module_cache_ram_248__7), .A1 (
             nx35636), .S0 (nx34516)) ;
    oai21 ix32906 (.Y (nx32905), .A0 (nx23880), .A1 (nx23802), .B0 (nx37268)) ;
    nand04 ix23881 (.Y (nx23880), .A0 (nx32908), .A1 (nx32916), .A2 (nx32924), .A3 (
           nx32932)) ;
    aoi22 ix32909 (.Y (nx32908), .A0 (camera_module_cache_ram_9__7), .A1 (
          nx35842), .B0 (camera_module_cache_ram_25__7), .B1 (nx35882)) ;
    dffr camera_module_cache_reg_ram_9__7 (.Q (camera_module_cache_ram_9__7), .QB (
         \$dummy [1966]), .D (nx20363), .CLK (clk), .R (rst)) ;
    mux21_ni ix20364 (.Y (nx20363), .A0 (camera_module_cache_ram_9__7), .A1 (
             nx35636), .S0 (nx34506)) ;
    dffr camera_module_cache_reg_ram_25__7 (.Q (camera_module_cache_ram_25__7), 
         .QB (\$dummy [1967]), .D (nx20353), .CLK (clk), .R (rst)) ;
    mux21_ni ix20354 (.Y (nx20353), .A0 (camera_module_cache_ram_25__7), .A1 (
             nx35636), .S0 (nx34502)) ;
    aoi22 ix32917 (.Y (nx32916), .A0 (camera_module_cache_ram_41__7), .A1 (
          nx35922), .B0 (camera_module_cache_ram_57__7), .B1 (nx35962)) ;
    dffr camera_module_cache_reg_ram_41__7 (.Q (camera_module_cache_ram_41__7), 
         .QB (\$dummy [1968]), .D (nx20343), .CLK (clk), .R (rst)) ;
    mux21_ni ix20344 (.Y (nx20343), .A0 (camera_module_cache_ram_41__7), .A1 (
             nx35636), .S0 (nx34498)) ;
    dffr camera_module_cache_reg_ram_57__7 (.Q (camera_module_cache_ram_57__7), 
         .QB (\$dummy [1969]), .D (nx20333), .CLK (clk), .R (rst)) ;
    mux21_ni ix20334 (.Y (nx20333), .A0 (camera_module_cache_ram_57__7), .A1 (
             nx35638), .S0 (nx34494)) ;
    aoi22 ix32925 (.Y (nx32924), .A0 (camera_module_cache_ram_73__7), .A1 (
          nx36002), .B0 (camera_module_cache_ram_89__7), .B1 (nx36042)) ;
    dffr camera_module_cache_reg_ram_73__7 (.Q (camera_module_cache_ram_73__7), 
         .QB (\$dummy [1970]), .D (nx20323), .CLK (clk), .R (rst)) ;
    mux21_ni ix20324 (.Y (nx20323), .A0 (camera_module_cache_ram_73__7), .A1 (
             nx35638), .S0 (nx34490)) ;
    dffr camera_module_cache_reg_ram_89__7 (.Q (camera_module_cache_ram_89__7), 
         .QB (\$dummy [1971]), .D (nx20313), .CLK (clk), .R (rst)) ;
    mux21_ni ix20314 (.Y (nx20313), .A0 (camera_module_cache_ram_89__7), .A1 (
             nx35638), .S0 (nx34486)) ;
    aoi22 ix32933 (.Y (nx32932), .A0 (camera_module_cache_ram_121__7), .A1 (
          nx36082), .B0 (camera_module_cache_ram_105__7), .B1 (nx36122)) ;
    dffr camera_module_cache_reg_ram_121__7 (.Q (camera_module_cache_ram_121__7)
         , .QB (\$dummy [1972]), .D (nx20293), .CLK (clk), .R (rst)) ;
    mux21_ni ix20294 (.Y (nx20293), .A0 (camera_module_cache_ram_121__7), .A1 (
             nx35638), .S0 (nx34478)) ;
    dffr camera_module_cache_reg_ram_105__7 (.Q (camera_module_cache_ram_105__7)
         , .QB (\$dummy [1973]), .D (nx20303), .CLK (clk), .R (rst)) ;
    mux21_ni ix20304 (.Y (nx20303), .A0 (camera_module_cache_ram_105__7), .A1 (
             nx35638), .S0 (nx34482)) ;
    nand04 ix23803 (.Y (nx23802), .A0 (nx32941), .A1 (nx32949), .A2 (nx32957), .A3 (
           nx32965)) ;
    aoi22 ix32942 (.Y (nx32941), .A0 (camera_module_cache_ram_137__7), .A1 (
          nx36162), .B0 (camera_module_cache_ram_153__7), .B1 (nx36202)) ;
    dffr camera_module_cache_reg_ram_137__7 (.Q (camera_module_cache_ram_137__7)
         , .QB (\$dummy [1974]), .D (nx20283), .CLK (clk), .R (rst)) ;
    mux21_ni ix20284 (.Y (nx20283), .A0 (camera_module_cache_ram_137__7), .A1 (
             nx35638), .S0 (nx34474)) ;
    dffr camera_module_cache_reg_ram_153__7 (.Q (camera_module_cache_ram_153__7)
         , .QB (\$dummy [1975]), .D (nx20273), .CLK (clk), .R (rst)) ;
    mux21_ni ix20274 (.Y (nx20273), .A0 (camera_module_cache_ram_153__7), .A1 (
             nx35638), .S0 (nx34470)) ;
    aoi22 ix32950 (.Y (nx32949), .A0 (camera_module_cache_ram_185__7), .A1 (
          nx36242), .B0 (camera_module_cache_ram_169__7), .B1 (nx36282)) ;
    dffr camera_module_cache_reg_ram_185__7 (.Q (camera_module_cache_ram_185__7)
         , .QB (\$dummy [1976]), .D (nx20253), .CLK (clk), .R (rst)) ;
    mux21_ni ix20254 (.Y (nx20253), .A0 (camera_module_cache_ram_185__7), .A1 (
             nx35640), .S0 (nx34462)) ;
    dffr camera_module_cache_reg_ram_169__7 (.Q (camera_module_cache_ram_169__7)
         , .QB (\$dummy [1977]), .D (nx20263), .CLK (clk), .R (rst)) ;
    mux21_ni ix20264 (.Y (nx20263), .A0 (camera_module_cache_ram_169__7), .A1 (
             nx35640), .S0 (nx34466)) ;
    aoi22 ix32958 (.Y (nx32957), .A0 (camera_module_cache_ram_201__7), .A1 (
          nx36322), .B0 (camera_module_cache_ram_217__7), .B1 (nx36362)) ;
    dffr camera_module_cache_reg_ram_201__7 (.Q (camera_module_cache_ram_201__7)
         , .QB (\$dummy [1978]), .D (nx20243), .CLK (clk), .R (rst)) ;
    mux21_ni ix20244 (.Y (nx20243), .A0 (camera_module_cache_ram_201__7), .A1 (
             nx35640), .S0 (nx34458)) ;
    dffr camera_module_cache_reg_ram_217__7 (.Q (camera_module_cache_ram_217__7)
         , .QB (\$dummy [1979]), .D (nx20233), .CLK (clk), .R (rst)) ;
    mux21_ni ix20234 (.Y (nx20233), .A0 (camera_module_cache_ram_217__7), .A1 (
             nx35640), .S0 (nx34454)) ;
    aoi22 ix32966 (.Y (nx32965), .A0 (camera_module_cache_ram_233__7), .A1 (
          nx36402), .B0 (camera_module_cache_ram_249__7), .B1 (nx36442)) ;
    dffr camera_module_cache_reg_ram_233__7 (.Q (camera_module_cache_ram_233__7)
         , .QB (\$dummy [1980]), .D (nx20223), .CLK (clk), .R (rst)) ;
    mux21_ni ix20224 (.Y (nx20223), .A0 (camera_module_cache_ram_233__7), .A1 (
             nx35640), .S0 (nx34450)) ;
    dffr camera_module_cache_reg_ram_249__7 (.Q (camera_module_cache_ram_249__7)
         , .QB (\$dummy [1981]), .D (nx20213), .CLK (clk), .R (rst)) ;
    mux21_ni ix20214 (.Y (nx20213), .A0 (camera_module_cache_ram_249__7), .A1 (
             nx35640), .S0 (nx34446)) ;
    oai21 ix32974 (.Y (nx32973), .A0 (nx23716), .A1 (nx23638), .B0 (nx37272)) ;
    nand04 ix23717 (.Y (nx23716), .A0 (nx32976), .A1 (nx32984), .A2 (nx32992), .A3 (
           nx33000)) ;
    aoi22 ix32977 (.Y (nx32976), .A0 (camera_module_cache_ram_10__7), .A1 (
          nx37200), .B0 (camera_module_cache_ram_26__7), .B1 (nx37202)) ;
    dffr camera_module_cache_reg_ram_10__7 (.Q (camera_module_cache_ram_10__7), 
         .QB (\$dummy [1982]), .D (nx20203), .CLK (clk), .R (rst)) ;
    mux21_ni ix20204 (.Y (nx20203), .A0 (camera_module_cache_ram_10__7), .A1 (
             nx35640), .S0 (nx34436)) ;
    dffr camera_module_cache_reg_ram_26__7 (.Q (camera_module_cache_ram_26__7), 
         .QB (\$dummy [1983]), .D (nx20193), .CLK (clk), .R (rst)) ;
    mux21_ni ix20194 (.Y (nx20193), .A0 (camera_module_cache_ram_26__7), .A1 (
             nx35642), .S0 (nx34432)) ;
    aoi22 ix32985 (.Y (nx32984), .A0 (camera_module_cache_ram_42__7), .A1 (
          nx37204), .B0 (camera_module_cache_ram_58__7), .B1 (nx37206)) ;
    dffr camera_module_cache_reg_ram_42__7 (.Q (camera_module_cache_ram_42__7), 
         .QB (\$dummy [1984]), .D (nx20183), .CLK (clk), .R (rst)) ;
    mux21_ni ix20184 (.Y (nx20183), .A0 (camera_module_cache_ram_42__7), .A1 (
             nx35642), .S0 (nx34428)) ;
    dffr camera_module_cache_reg_ram_58__7 (.Q (camera_module_cache_ram_58__7), 
         .QB (\$dummy [1985]), .D (nx20173), .CLK (clk), .R (rst)) ;
    mux21_ni ix20174 (.Y (nx20173), .A0 (camera_module_cache_ram_58__7), .A1 (
             nx35642), .S0 (nx34424)) ;
    aoi22 ix32993 (.Y (nx32992), .A0 (camera_module_cache_ram_74__7), .A1 (
          nx37208), .B0 (camera_module_cache_ram_90__7), .B1 (nx37210)) ;
    dffr camera_module_cache_reg_ram_74__7 (.Q (camera_module_cache_ram_74__7), 
         .QB (\$dummy [1986]), .D (nx20163), .CLK (clk), .R (rst)) ;
    mux21_ni ix20164 (.Y (nx20163), .A0 (camera_module_cache_ram_74__7), .A1 (
             nx35642), .S0 (nx34420)) ;
    dffr camera_module_cache_reg_ram_90__7 (.Q (camera_module_cache_ram_90__7), 
         .QB (\$dummy [1987]), .D (nx20153), .CLK (clk), .R (rst)) ;
    mux21_ni ix20154 (.Y (nx20153), .A0 (camera_module_cache_ram_90__7), .A1 (
             nx35642), .S0 (nx34416)) ;
    aoi22 ix33001 (.Y (nx33000), .A0 (camera_module_cache_ram_122__7), .A1 (
          nx37212), .B0 (camera_module_cache_ram_106__7), .B1 (nx37214)) ;
    dffr camera_module_cache_reg_ram_122__7 (.Q (camera_module_cache_ram_122__7)
         , .QB (\$dummy [1988]), .D (nx20133), .CLK (clk), .R (rst)) ;
    mux21_ni ix20134 (.Y (nx20133), .A0 (camera_module_cache_ram_122__7), .A1 (
             nx35642), .S0 (nx34408)) ;
    dffr camera_module_cache_reg_ram_106__7 (.Q (camera_module_cache_ram_106__7)
         , .QB (\$dummy [1989]), .D (nx20143), .CLK (clk), .R (rst)) ;
    mux21_ni ix20144 (.Y (nx20143), .A0 (camera_module_cache_ram_106__7), .A1 (
             nx35642), .S0 (nx34412)) ;
    nand04 ix23639 (.Y (nx23638), .A0 (nx33009), .A1 (nx33017), .A2 (nx33025), .A3 (
           nx33033)) ;
    aoi22 ix33010 (.Y (nx33009), .A0 (camera_module_cache_ram_138__7), .A1 (
          nx37216), .B0 (camera_module_cache_ram_154__7), .B1 (nx37218)) ;
    dffr camera_module_cache_reg_ram_138__7 (.Q (camera_module_cache_ram_138__7)
         , .QB (\$dummy [1990]), .D (nx20123), .CLK (clk), .R (rst)) ;
    mux21_ni ix20124 (.Y (nx20123), .A0 (camera_module_cache_ram_138__7), .A1 (
             nx35644), .S0 (nx34404)) ;
    dffr camera_module_cache_reg_ram_154__7 (.Q (camera_module_cache_ram_154__7)
         , .QB (\$dummy [1991]), .D (nx20113), .CLK (clk), .R (rst)) ;
    mux21_ni ix20114 (.Y (nx20113), .A0 (camera_module_cache_ram_154__7), .A1 (
             nx35644), .S0 (nx34400)) ;
    aoi22 ix33018 (.Y (nx33017), .A0 (camera_module_cache_ram_186__7), .A1 (
          nx37220), .B0 (camera_module_cache_ram_170__7), .B1 (nx37222)) ;
    dffr camera_module_cache_reg_ram_186__7 (.Q (camera_module_cache_ram_186__7)
         , .QB (\$dummy [1992]), .D (nx20093), .CLK (clk), .R (rst)) ;
    mux21_ni ix20094 (.Y (nx20093), .A0 (camera_module_cache_ram_186__7), .A1 (
             nx35644), .S0 (nx34392)) ;
    dffr camera_module_cache_reg_ram_170__7 (.Q (camera_module_cache_ram_170__7)
         , .QB (\$dummy [1993]), .D (nx20103), .CLK (clk), .R (rst)) ;
    mux21_ni ix20104 (.Y (nx20103), .A0 (camera_module_cache_ram_170__7), .A1 (
             nx35644), .S0 (nx34396)) ;
    aoi22 ix33026 (.Y (nx33025), .A0 (camera_module_cache_ram_202__7), .A1 (
          nx37224), .B0 (camera_module_cache_ram_218__7), .B1 (nx37226)) ;
    dffr camera_module_cache_reg_ram_202__7 (.Q (camera_module_cache_ram_202__7)
         , .QB (\$dummy [1994]), .D (nx20083), .CLK (clk), .R (rst)) ;
    mux21_ni ix20084 (.Y (nx20083), .A0 (camera_module_cache_ram_202__7), .A1 (
             nx35644), .S0 (nx34388)) ;
    dffr camera_module_cache_reg_ram_218__7 (.Q (camera_module_cache_ram_218__7)
         , .QB (\$dummy [1995]), .D (nx20073), .CLK (clk), .R (rst)) ;
    mux21_ni ix20074 (.Y (nx20073), .A0 (camera_module_cache_ram_218__7), .A1 (
             nx35644), .S0 (nx34384)) ;
    aoi22 ix33034 (.Y (nx33033), .A0 (camera_module_cache_ram_234__7), .A1 (
          nx37228), .B0 (camera_module_cache_ram_250__7), .B1 (nx37230)) ;
    dffr camera_module_cache_reg_ram_234__7 (.Q (camera_module_cache_ram_234__7)
         , .QB (\$dummy [1996]), .D (nx20063), .CLK (clk), .R (rst)) ;
    mux21_ni ix20064 (.Y (nx20063), .A0 (camera_module_cache_ram_234__7), .A1 (
             nx35644), .S0 (nx34380)) ;
    dffr camera_module_cache_reg_ram_250__7 (.Q (camera_module_cache_ram_250__7)
         , .QB (\$dummy [1997]), .D (nx20053), .CLK (clk), .R (rst)) ;
    mux21_ni ix20054 (.Y (nx20053), .A0 (camera_module_cache_ram_250__7), .A1 (
             nx35646), .S0 (nx34376)) ;
    oai21 ix33042 (.Y (nx33041), .A0 (nx23554), .A1 (nx23476), .B0 (nx37276)) ;
    nand04 ix23555 (.Y (nx23554), .A0 (nx33044), .A1 (nx33052), .A2 (nx33060), .A3 (
           nx33068)) ;
    aoi22 ix33045 (.Y (nx33044), .A0 (camera_module_cache_ram_11__7), .A1 (
          nx37200), .B0 (camera_module_cache_ram_27__7), .B1 (nx37202)) ;
    dffr camera_module_cache_reg_ram_11__7 (.Q (camera_module_cache_ram_11__7), 
         .QB (\$dummy [1998]), .D (nx20043), .CLK (clk), .R (rst)) ;
    mux21_ni ix20044 (.Y (nx20043), .A0 (camera_module_cache_ram_11__7), .A1 (
             nx35646), .S0 (nx34366)) ;
    dffr camera_module_cache_reg_ram_27__7 (.Q (camera_module_cache_ram_27__7), 
         .QB (\$dummy [1999]), .D (nx20033), .CLK (clk), .R (rst)) ;
    mux21_ni ix20034 (.Y (nx20033), .A0 (camera_module_cache_ram_27__7), .A1 (
             nx35646), .S0 (nx34362)) ;
    aoi22 ix33053 (.Y (nx33052), .A0 (camera_module_cache_ram_43__7), .A1 (
          nx37204), .B0 (camera_module_cache_ram_59__7), .B1 (nx37206)) ;
    dffr camera_module_cache_reg_ram_43__7 (.Q (camera_module_cache_ram_43__7), 
         .QB (\$dummy [2000]), .D (nx20023), .CLK (clk), .R (rst)) ;
    mux21_ni ix20024 (.Y (nx20023), .A0 (camera_module_cache_ram_43__7), .A1 (
             nx35646), .S0 (nx34358)) ;
    dffr camera_module_cache_reg_ram_59__7 (.Q (camera_module_cache_ram_59__7), 
         .QB (\$dummy [2001]), .D (nx20013), .CLK (clk), .R (rst)) ;
    mux21_ni ix20014 (.Y (nx20013), .A0 (camera_module_cache_ram_59__7), .A1 (
             nx35646), .S0 (nx34354)) ;
    aoi22 ix33061 (.Y (nx33060), .A0 (camera_module_cache_ram_75__7), .A1 (
          nx37208), .B0 (camera_module_cache_ram_91__7), .B1 (nx37210)) ;
    dffr camera_module_cache_reg_ram_75__7 (.Q (camera_module_cache_ram_75__7), 
         .QB (\$dummy [2002]), .D (nx20003), .CLK (clk), .R (rst)) ;
    mux21_ni ix20004 (.Y (nx20003), .A0 (camera_module_cache_ram_75__7), .A1 (
             nx35646), .S0 (nx34350)) ;
    dffr camera_module_cache_reg_ram_91__7 (.Q (camera_module_cache_ram_91__7), 
         .QB (\$dummy [2003]), .D (nx19993), .CLK (clk), .R (rst)) ;
    mux21_ni ix19994 (.Y (nx19993), .A0 (camera_module_cache_ram_91__7), .A1 (
             nx35646), .S0 (nx34346)) ;
    aoi22 ix33069 (.Y (nx33068), .A0 (camera_module_cache_ram_123__7), .A1 (
          nx37212), .B0 (camera_module_cache_ram_107__7), .B1 (nx37214)) ;
    dffr camera_module_cache_reg_ram_123__7 (.Q (camera_module_cache_ram_123__7)
         , .QB (\$dummy [2004]), .D (nx19973), .CLK (clk), .R (rst)) ;
    mux21_ni ix19974 (.Y (nx19973), .A0 (camera_module_cache_ram_123__7), .A1 (
             nx35648), .S0 (nx34338)) ;
    dffr camera_module_cache_reg_ram_107__7 (.Q (camera_module_cache_ram_107__7)
         , .QB (\$dummy [2005]), .D (nx19983), .CLK (clk), .R (rst)) ;
    mux21_ni ix19984 (.Y (nx19983), .A0 (camera_module_cache_ram_107__7), .A1 (
             nx35648), .S0 (nx34342)) ;
    nand04 ix23477 (.Y (nx23476), .A0 (nx33077), .A1 (nx33085), .A2 (nx33093), .A3 (
           nx33101)) ;
    aoi22 ix33078 (.Y (nx33077), .A0 (camera_module_cache_ram_139__7), .A1 (
          nx37216), .B0 (camera_module_cache_ram_155__7), .B1 (nx37218)) ;
    dffr camera_module_cache_reg_ram_139__7 (.Q (camera_module_cache_ram_139__7)
         , .QB (\$dummy [2006]), .D (nx19963), .CLK (clk), .R (rst)) ;
    mux21_ni ix19964 (.Y (nx19963), .A0 (camera_module_cache_ram_139__7), .A1 (
             nx35648), .S0 (nx34334)) ;
    dffr camera_module_cache_reg_ram_155__7 (.Q (camera_module_cache_ram_155__7)
         , .QB (\$dummy [2007]), .D (nx19953), .CLK (clk), .R (rst)) ;
    mux21_ni ix19954 (.Y (nx19953), .A0 (camera_module_cache_ram_155__7), .A1 (
             nx35648), .S0 (nx34330)) ;
    aoi22 ix33086 (.Y (nx33085), .A0 (camera_module_cache_ram_187__7), .A1 (
          nx37220), .B0 (camera_module_cache_ram_171__7), .B1 (nx37222)) ;
    dffr camera_module_cache_reg_ram_187__7 (.Q (camera_module_cache_ram_187__7)
         , .QB (\$dummy [2008]), .D (nx19933), .CLK (clk), .R (rst)) ;
    mux21_ni ix19934 (.Y (nx19933), .A0 (camera_module_cache_ram_187__7), .A1 (
             nx35648), .S0 (nx34322)) ;
    dffr camera_module_cache_reg_ram_171__7 (.Q (camera_module_cache_ram_171__7)
         , .QB (\$dummy [2009]), .D (nx19943), .CLK (clk), .R (rst)) ;
    mux21_ni ix19944 (.Y (nx19943), .A0 (camera_module_cache_ram_171__7), .A1 (
             nx35648), .S0 (nx34326)) ;
    aoi22 ix33094 (.Y (nx33093), .A0 (camera_module_cache_ram_203__7), .A1 (
          nx37224), .B0 (camera_module_cache_ram_219__7), .B1 (nx37226)) ;
    dffr camera_module_cache_reg_ram_203__7 (.Q (camera_module_cache_ram_203__7)
         , .QB (\$dummy [2010]), .D (nx19923), .CLK (clk), .R (rst)) ;
    mux21_ni ix19924 (.Y (nx19923), .A0 (camera_module_cache_ram_203__7), .A1 (
             nx35648), .S0 (nx34318)) ;
    dffr camera_module_cache_reg_ram_219__7 (.Q (camera_module_cache_ram_219__7)
         , .QB (\$dummy [2011]), .D (nx19913), .CLK (clk), .R (rst)) ;
    mux21_ni ix19914 (.Y (nx19913), .A0 (camera_module_cache_ram_219__7), .A1 (
             nx35650), .S0 (nx34314)) ;
    aoi22 ix33102 (.Y (nx33101), .A0 (camera_module_cache_ram_235__7), .A1 (
          nx37228), .B0 (camera_module_cache_ram_251__7), .B1 (nx37230)) ;
    dffr camera_module_cache_reg_ram_235__7 (.Q (camera_module_cache_ram_235__7)
         , .QB (\$dummy [2012]), .D (nx19903), .CLK (clk), .R (rst)) ;
    mux21_ni ix19904 (.Y (nx19903), .A0 (camera_module_cache_ram_235__7), .A1 (
             nx35650), .S0 (nx34310)) ;
    dffr camera_module_cache_reg_ram_251__7 (.Q (camera_module_cache_ram_251__7)
         , .QB (\$dummy [2013]), .D (nx19893), .CLK (clk), .R (rst)) ;
    mux21_ni ix19894 (.Y (nx19893), .A0 (camera_module_cache_ram_251__7), .A1 (
             nx35650), .S0 (nx34306)) ;
    nand04 ix23399 (.Y (nx23398), .A0 (nx33110), .A1 (nx33178), .A2 (nx33246), .A3 (
           nx33314)) ;
    oai21 ix33111 (.Y (nx33110), .A0 (nx23388), .A1 (nx23310), .B0 (nx36508)) ;
    nand04 ix23389 (.Y (nx23388), .A0 (nx33113), .A1 (nx33121), .A2 (nx33129), .A3 (
           nx33137)) ;
    aoi22 ix33114 (.Y (nx33113), .A0 (camera_module_cache_ram_12__7), .A1 (
          nx37200), .B0 (camera_module_cache_ram_28__7), .B1 (nx37202)) ;
    dffr camera_module_cache_reg_ram_12__7 (.Q (camera_module_cache_ram_12__7), 
         .QB (\$dummy [2014]), .D (nx19883), .CLK (clk), .R (rst)) ;
    mux21_ni ix19884 (.Y (nx19883), .A0 (nx35650), .A1 (
             camera_module_cache_ram_12__7), .S0 (nx36498)) ;
    dffr camera_module_cache_reg_ram_28__7 (.Q (camera_module_cache_ram_28__7), 
         .QB (\$dummy [2015]), .D (nx19873), .CLK (clk), .R (rst)) ;
    mux21_ni ix19874 (.Y (nx19873), .A0 (nx35650), .A1 (
             camera_module_cache_ram_28__7), .S0 (nx36512)) ;
    aoi22 ix33122 (.Y (nx33121), .A0 (camera_module_cache_ram_44__7), .A1 (
          nx37204), .B0 (camera_module_cache_ram_60__7), .B1 (nx37206)) ;
    dffr camera_module_cache_reg_ram_44__7 (.Q (camera_module_cache_ram_44__7), 
         .QB (\$dummy [2016]), .D (nx19863), .CLK (clk), .R (rst)) ;
    mux21_ni ix19864 (.Y (nx19863), .A0 (nx35650), .A1 (
             camera_module_cache_ram_44__7), .S0 (nx36516)) ;
    dffr camera_module_cache_reg_ram_60__7 (.Q (camera_module_cache_ram_60__7), 
         .QB (\$dummy [2017]), .D (nx19853), .CLK (clk), .R (rst)) ;
    mux21_ni ix19854 (.Y (nx19853), .A0 (nx35650), .A1 (
             camera_module_cache_ram_60__7), .S0 (nx36520)) ;
    aoi22 ix33130 (.Y (nx33129), .A0 (camera_module_cache_ram_76__7), .A1 (
          nx37208), .B0 (camera_module_cache_ram_92__7), .B1 (nx37210)) ;
    dffr camera_module_cache_reg_ram_76__7 (.Q (camera_module_cache_ram_76__7), 
         .QB (\$dummy [2018]), .D (nx19843), .CLK (clk), .R (rst)) ;
    mux21_ni ix19844 (.Y (nx19843), .A0 (nx35652), .A1 (
             camera_module_cache_ram_76__7), .S0 (nx36524)) ;
    dffr camera_module_cache_reg_ram_92__7 (.Q (camera_module_cache_ram_92__7), 
         .QB (\$dummy [2019]), .D (nx19833), .CLK (clk), .R (rst)) ;
    mux21_ni ix19834 (.Y (nx19833), .A0 (nx35652), .A1 (
             camera_module_cache_ram_92__7), .S0 (nx36528)) ;
    aoi22 ix33138 (.Y (nx33137), .A0 (camera_module_cache_ram_124__7), .A1 (
          nx37212), .B0 (camera_module_cache_ram_108__7), .B1 (nx37214)) ;
    dffr camera_module_cache_reg_ram_124__7 (.Q (camera_module_cache_ram_124__7)
         , .QB (\$dummy [2020]), .D (nx19813), .CLK (clk), .R (rst)) ;
    mux21_ni ix19814 (.Y (nx19813), .A0 (nx35652), .A1 (
             camera_module_cache_ram_124__7), .S0 (nx36532)) ;
    dffr camera_module_cache_reg_ram_108__7 (.Q (camera_module_cache_ram_108__7)
         , .QB (\$dummy [2021]), .D (nx19823), .CLK (clk), .R (rst)) ;
    mux21_ni ix19824 (.Y (nx19823), .A0 (nx35652), .A1 (
             camera_module_cache_ram_108__7), .S0 (nx36536)) ;
    nand04 ix23311 (.Y (nx23310), .A0 (nx33146), .A1 (nx33154), .A2 (nx33162), .A3 (
           nx33170)) ;
    aoi22 ix33147 (.Y (nx33146), .A0 (camera_module_cache_ram_140__7), .A1 (
          nx37216), .B0 (camera_module_cache_ram_156__7), .B1 (nx37218)) ;
    dffr camera_module_cache_reg_ram_140__7 (.Q (camera_module_cache_ram_140__7)
         , .QB (\$dummy [2022]), .D (nx19803), .CLK (clk), .R (rst)) ;
    mux21_ni ix19804 (.Y (nx19803), .A0 (nx35652), .A1 (
             camera_module_cache_ram_140__7), .S0 (nx36540)) ;
    dffr camera_module_cache_reg_ram_156__7 (.Q (camera_module_cache_ram_156__7)
         , .QB (\$dummy [2023]), .D (nx19793), .CLK (clk), .R (rst)) ;
    mux21_ni ix19794 (.Y (nx19793), .A0 (nx35652), .A1 (
             camera_module_cache_ram_156__7), .S0 (nx36544)) ;
    aoi22 ix33155 (.Y (nx33154), .A0 (camera_module_cache_ram_188__7), .A1 (
          nx37220), .B0 (camera_module_cache_ram_172__7), .B1 (nx37222)) ;
    dffr camera_module_cache_reg_ram_188__7 (.Q (camera_module_cache_ram_188__7)
         , .QB (\$dummy [2024]), .D (nx19773), .CLK (clk), .R (rst)) ;
    mux21_ni ix19774 (.Y (nx19773), .A0 (nx35652), .A1 (
             camera_module_cache_ram_188__7), .S0 (nx36548)) ;
    dffr camera_module_cache_reg_ram_172__7 (.Q (camera_module_cache_ram_172__7)
         , .QB (\$dummy [2025]), .D (nx19783), .CLK (clk), .R (rst)) ;
    mux21_ni ix19784 (.Y (nx19783), .A0 (nx35654), .A1 (
             camera_module_cache_ram_172__7), .S0 (nx36552)) ;
    aoi22 ix33163 (.Y (nx33162), .A0 (camera_module_cache_ram_204__7), .A1 (
          nx37224), .B0 (camera_module_cache_ram_220__7), .B1 (nx37226)) ;
    dffr camera_module_cache_reg_ram_204__7 (.Q (camera_module_cache_ram_204__7)
         , .QB (\$dummy [2026]), .D (nx19763), .CLK (clk), .R (rst)) ;
    mux21_ni ix19764 (.Y (nx19763), .A0 (nx35654), .A1 (
             camera_module_cache_ram_204__7), .S0 (nx36556)) ;
    dffr camera_module_cache_reg_ram_220__7 (.Q (camera_module_cache_ram_220__7)
         , .QB (\$dummy [2027]), .D (nx19753), .CLK (clk), .R (rst)) ;
    mux21_ni ix19754 (.Y (nx19753), .A0 (nx35654), .A1 (
             camera_module_cache_ram_220__7), .S0 (nx36560)) ;
    aoi22 ix33171 (.Y (nx33170), .A0 (camera_module_cache_ram_236__7), .A1 (
          nx37228), .B0 (camera_module_cache_ram_252__7), .B1 (nx37230)) ;
    dffr camera_module_cache_reg_ram_236__7 (.Q (camera_module_cache_ram_236__7)
         , .QB (\$dummy [2028]), .D (nx19743), .CLK (clk), .R (rst)) ;
    mux21_ni ix19744 (.Y (nx19743), .A0 (nx35654), .A1 (
             camera_module_cache_ram_236__7), .S0 (nx36564)) ;
    dffr camera_module_cache_reg_ram_252__7 (.Q (camera_module_cache_ram_252__7)
         , .QB (\$dummy [2029]), .D (nx19733), .CLK (clk), .R (rst)) ;
    mux21_ni ix19734 (.Y (nx19733), .A0 (nx35654), .A1 (
             camera_module_cache_ram_252__7), .S0 (nx36568)) ;
    oai21 ix33179 (.Y (nx33178), .A0 (nx23226), .A1 (nx23148), .B0 (nx36582)) ;
    nand04 ix23227 (.Y (nx23226), .A0 (nx33181), .A1 (nx33189), .A2 (nx33197), .A3 (
           nx33205)) ;
    aoi22 ix33182 (.Y (nx33181), .A0 (camera_module_cache_ram_13__7), .A1 (
          nx37200), .B0 (camera_module_cache_ram_29__7), .B1 (nx37202)) ;
    dffr camera_module_cache_reg_ram_13__7 (.Q (camera_module_cache_ram_13__7), 
         .QB (\$dummy [2030]), .D (nx19723), .CLK (clk), .R (rst)) ;
    mux21_ni ix19724 (.Y (nx19723), .A0 (nx35654), .A1 (
             camera_module_cache_ram_13__7), .S0 (nx36572)) ;
    dffr camera_module_cache_reg_ram_29__7 (.Q (camera_module_cache_ram_29__7), 
         .QB (\$dummy [2031]), .D (nx19713), .CLK (clk), .R (rst)) ;
    mux21_ni ix19714 (.Y (nx19713), .A0 (nx35654), .A1 (
             camera_module_cache_ram_29__7), .S0 (nx36586)) ;
    aoi22 ix33190 (.Y (nx33189), .A0 (camera_module_cache_ram_45__7), .A1 (
          nx37204), .B0 (camera_module_cache_ram_61__7), .B1 (nx37206)) ;
    dffr camera_module_cache_reg_ram_45__7 (.Q (camera_module_cache_ram_45__7), 
         .QB (\$dummy [2032]), .D (nx19703), .CLK (clk), .R (rst)) ;
    mux21_ni ix19704 (.Y (nx19703), .A0 (nx35656), .A1 (
             camera_module_cache_ram_45__7), .S0 (nx36590)) ;
    dffr camera_module_cache_reg_ram_61__7 (.Q (camera_module_cache_ram_61__7), 
         .QB (\$dummy [2033]), .D (nx19693), .CLK (clk), .R (rst)) ;
    mux21_ni ix19694 (.Y (nx19693), .A0 (nx35656), .A1 (
             camera_module_cache_ram_61__7), .S0 (nx36594)) ;
    aoi22 ix33198 (.Y (nx33197), .A0 (camera_module_cache_ram_77__7), .A1 (
          nx37208), .B0 (camera_module_cache_ram_93__7), .B1 (nx37210)) ;
    dffr camera_module_cache_reg_ram_77__7 (.Q (camera_module_cache_ram_77__7), 
         .QB (\$dummy [2034]), .D (nx19683), .CLK (clk), .R (rst)) ;
    mux21_ni ix19684 (.Y (nx19683), .A0 (nx35656), .A1 (
             camera_module_cache_ram_77__7), .S0 (nx36598)) ;
    dffr camera_module_cache_reg_ram_93__7 (.Q (camera_module_cache_ram_93__7), 
         .QB (\$dummy [2035]), .D (nx19673), .CLK (clk), .R (rst)) ;
    mux21_ni ix19674 (.Y (nx19673), .A0 (nx35656), .A1 (
             camera_module_cache_ram_93__7), .S0 (nx36602)) ;
    aoi22 ix33206 (.Y (nx33205), .A0 (camera_module_cache_ram_125__7), .A1 (
          nx37212), .B0 (camera_module_cache_ram_109__7), .B1 (nx37214)) ;
    dffr camera_module_cache_reg_ram_125__7 (.Q (camera_module_cache_ram_125__7)
         , .QB (\$dummy [2036]), .D (nx19653), .CLK (clk), .R (rst)) ;
    mux21_ni ix19654 (.Y (nx19653), .A0 (nx35656), .A1 (
             camera_module_cache_ram_125__7), .S0 (nx36606)) ;
    dffr camera_module_cache_reg_ram_109__7 (.Q (camera_module_cache_ram_109__7)
         , .QB (\$dummy [2037]), .D (nx19663), .CLK (clk), .R (rst)) ;
    mux21_ni ix19664 (.Y (nx19663), .A0 (nx35656), .A1 (
             camera_module_cache_ram_109__7), .S0 (nx36610)) ;
    nand04 ix23149 (.Y (nx23148), .A0 (nx33214), .A1 (nx33222), .A2 (nx33230), .A3 (
           nx33238)) ;
    aoi22 ix33215 (.Y (nx33214), .A0 (camera_module_cache_ram_141__7), .A1 (
          nx37216), .B0 (camera_module_cache_ram_157__7), .B1 (nx37218)) ;
    dffr camera_module_cache_reg_ram_141__7 (.Q (camera_module_cache_ram_141__7)
         , .QB (\$dummy [2038]), .D (nx19643), .CLK (clk), .R (rst)) ;
    mux21_ni ix19644 (.Y (nx19643), .A0 (nx35656), .A1 (
             camera_module_cache_ram_141__7), .S0 (nx36614)) ;
    dffr camera_module_cache_reg_ram_157__7 (.Q (camera_module_cache_ram_157__7)
         , .QB (\$dummy [2039]), .D (nx19633), .CLK (clk), .R (rst)) ;
    mux21_ni ix19634 (.Y (nx19633), .A0 (nx35658), .A1 (
             camera_module_cache_ram_157__7), .S0 (nx36618)) ;
    aoi22 ix33223 (.Y (nx33222), .A0 (camera_module_cache_ram_189__7), .A1 (
          nx37220), .B0 (camera_module_cache_ram_173__7), .B1 (nx37222)) ;
    dffr camera_module_cache_reg_ram_189__7 (.Q (camera_module_cache_ram_189__7)
         , .QB (\$dummy [2040]), .D (nx19613), .CLK (clk), .R (rst)) ;
    mux21_ni ix19614 (.Y (nx19613), .A0 (nx35658), .A1 (
             camera_module_cache_ram_189__7), .S0 (nx36622)) ;
    dffr camera_module_cache_reg_ram_173__7 (.Q (camera_module_cache_ram_173__7)
         , .QB (\$dummy [2041]), .D (nx19623), .CLK (clk), .R (rst)) ;
    mux21_ni ix19624 (.Y (nx19623), .A0 (nx35658), .A1 (
             camera_module_cache_ram_173__7), .S0 (nx36626)) ;
    aoi22 ix33231 (.Y (nx33230), .A0 (camera_module_cache_ram_205__7), .A1 (
          nx37224), .B0 (camera_module_cache_ram_221__7), .B1 (nx37226)) ;
    dffr camera_module_cache_reg_ram_205__7 (.Q (camera_module_cache_ram_205__7)
         , .QB (\$dummy [2042]), .D (nx19603), .CLK (clk), .R (rst)) ;
    mux21_ni ix19604 (.Y (nx19603), .A0 (nx35658), .A1 (
             camera_module_cache_ram_205__7), .S0 (nx36630)) ;
    dffr camera_module_cache_reg_ram_221__7 (.Q (camera_module_cache_ram_221__7)
         , .QB (\$dummy [2043]), .D (nx19593), .CLK (clk), .R (rst)) ;
    mux21_ni ix19594 (.Y (nx19593), .A0 (nx35658), .A1 (
             camera_module_cache_ram_221__7), .S0 (nx36634)) ;
    aoi22 ix33239 (.Y (nx33238), .A0 (camera_module_cache_ram_237__7), .A1 (
          nx37228), .B0 (camera_module_cache_ram_253__7), .B1 (nx37230)) ;
    dffr camera_module_cache_reg_ram_237__7 (.Q (camera_module_cache_ram_237__7)
         , .QB (\$dummy [2044]), .D (nx19583), .CLK (clk), .R (rst)) ;
    mux21_ni ix19584 (.Y (nx19583), .A0 (nx35658), .A1 (
             camera_module_cache_ram_237__7), .S0 (nx36638)) ;
    dffr camera_module_cache_reg_ram_253__7 (.Q (camera_module_cache_ram_253__7)
         , .QB (\$dummy [2045]), .D (nx19573), .CLK (clk), .R (rst)) ;
    mux21_ni ix19574 (.Y (nx19573), .A0 (nx35658), .A1 (
             camera_module_cache_ram_253__7), .S0 (nx36642)) ;
    oai21 ix33247 (.Y (nx33246), .A0 (nx23062), .A1 (nx22984), .B0 (nx36656)) ;
    nand04 ix23063 (.Y (nx23062), .A0 (nx33249), .A1 (nx33257), .A2 (nx33265), .A3 (
           nx33273)) ;
    aoi22 ix33250 (.Y (nx33249), .A0 (camera_module_cache_ram_14__7), .A1 (
          nx37200), .B0 (camera_module_cache_ram_30__7), .B1 (nx37202)) ;
    dffr camera_module_cache_reg_ram_14__7 (.Q (camera_module_cache_ram_14__7), 
         .QB (\$dummy [2046]), .D (nx19563), .CLK (clk), .R (rst)) ;
    mux21_ni ix19564 (.Y (nx19563), .A0 (nx35660), .A1 (
             camera_module_cache_ram_14__7), .S0 (nx36646)) ;
    dffr camera_module_cache_reg_ram_30__7 (.Q (camera_module_cache_ram_30__7), 
         .QB (\$dummy [2047]), .D (nx19553), .CLK (clk), .R (rst)) ;
    mux21_ni ix19554 (.Y (nx19553), .A0 (nx35660), .A1 (
             camera_module_cache_ram_30__7), .S0 (nx36660)) ;
    aoi22 ix33258 (.Y (nx33257), .A0 (camera_module_cache_ram_46__7), .A1 (
          nx37204), .B0 (camera_module_cache_ram_62__7), .B1 (nx37206)) ;
    dffr camera_module_cache_reg_ram_46__7 (.Q (camera_module_cache_ram_46__7), 
         .QB (\$dummy [2048]), .D (nx19543), .CLK (clk), .R (rst)) ;
    mux21_ni ix19544 (.Y (nx19543), .A0 (nx35660), .A1 (
             camera_module_cache_ram_46__7), .S0 (nx36664)) ;
    dffr camera_module_cache_reg_ram_62__7 (.Q (camera_module_cache_ram_62__7), 
         .QB (\$dummy [2049]), .D (nx19533), .CLK (clk), .R (rst)) ;
    mux21_ni ix19534 (.Y (nx19533), .A0 (nx35660), .A1 (
             camera_module_cache_ram_62__7), .S0 (nx36668)) ;
    aoi22 ix33266 (.Y (nx33265), .A0 (camera_module_cache_ram_78__7), .A1 (
          nx37208), .B0 (camera_module_cache_ram_94__7), .B1 (nx37210)) ;
    dffr camera_module_cache_reg_ram_78__7 (.Q (camera_module_cache_ram_78__7), 
         .QB (\$dummy [2050]), .D (nx19523), .CLK (clk), .R (rst)) ;
    mux21_ni ix19524 (.Y (nx19523), .A0 (nx35660), .A1 (
             camera_module_cache_ram_78__7), .S0 (nx36672)) ;
    dffr camera_module_cache_reg_ram_94__7 (.Q (camera_module_cache_ram_94__7), 
         .QB (\$dummy [2051]), .D (nx19513), .CLK (clk), .R (rst)) ;
    mux21_ni ix19514 (.Y (nx19513), .A0 (nx35660), .A1 (
             camera_module_cache_ram_94__7), .S0 (nx36676)) ;
    aoi22 ix33274 (.Y (nx33273), .A0 (camera_module_cache_ram_126__7), .A1 (
          nx37212), .B0 (camera_module_cache_ram_110__7), .B1 (nx37214)) ;
    dffr camera_module_cache_reg_ram_126__7 (.Q (camera_module_cache_ram_126__7)
         , .QB (\$dummy [2052]), .D (nx19493), .CLK (clk), .R (rst)) ;
    mux21_ni ix19494 (.Y (nx19493), .A0 (nx35660), .A1 (
             camera_module_cache_ram_126__7), .S0 (nx36680)) ;
    dffr camera_module_cache_reg_ram_110__7 (.Q (camera_module_cache_ram_110__7)
         , .QB (\$dummy [2053]), .D (nx19503), .CLK (clk), .R (rst)) ;
    mux21_ni ix19504 (.Y (nx19503), .A0 (nx35662), .A1 (
             camera_module_cache_ram_110__7), .S0 (nx36684)) ;
    nand04 ix22985 (.Y (nx22984), .A0 (nx33282), .A1 (nx33290), .A2 (nx33298), .A3 (
           nx33306)) ;
    aoi22 ix33283 (.Y (nx33282), .A0 (camera_module_cache_ram_142__7), .A1 (
          nx37216), .B0 (camera_module_cache_ram_158__7), .B1 (nx37218)) ;
    dffr camera_module_cache_reg_ram_142__7 (.Q (camera_module_cache_ram_142__7)
         , .QB (\$dummy [2054]), .D (nx19483), .CLK (clk), .R (rst)) ;
    mux21_ni ix19484 (.Y (nx19483), .A0 (nx35662), .A1 (
             camera_module_cache_ram_142__7), .S0 (nx36688)) ;
    dffr camera_module_cache_reg_ram_158__7 (.Q (camera_module_cache_ram_158__7)
         , .QB (\$dummy [2055]), .D (nx19473), .CLK (clk), .R (rst)) ;
    mux21_ni ix19474 (.Y (nx19473), .A0 (nx35662), .A1 (
             camera_module_cache_ram_158__7), .S0 (nx36692)) ;
    aoi22 ix33291 (.Y (nx33290), .A0 (camera_module_cache_ram_190__7), .A1 (
          nx37220), .B0 (camera_module_cache_ram_174__7), .B1 (nx37222)) ;
    dffr camera_module_cache_reg_ram_190__7 (.Q (camera_module_cache_ram_190__7)
         , .QB (\$dummy [2056]), .D (nx19453), .CLK (clk), .R (rst)) ;
    mux21_ni ix19454 (.Y (nx19453), .A0 (nx35662), .A1 (
             camera_module_cache_ram_190__7), .S0 (nx36696)) ;
    dffr camera_module_cache_reg_ram_174__7 (.Q (camera_module_cache_ram_174__7)
         , .QB (\$dummy [2057]), .D (nx19463), .CLK (clk), .R (rst)) ;
    mux21_ni ix19464 (.Y (nx19463), .A0 (nx35662), .A1 (
             camera_module_cache_ram_174__7), .S0 (nx36700)) ;
    aoi22 ix33299 (.Y (nx33298), .A0 (camera_module_cache_ram_206__7), .A1 (
          nx37224), .B0 (camera_module_cache_ram_222__7), .B1 (nx37226)) ;
    dffr camera_module_cache_reg_ram_206__7 (.Q (camera_module_cache_ram_206__7)
         , .QB (\$dummy [2058]), .D (nx19443), .CLK (clk), .R (rst)) ;
    mux21_ni ix19444 (.Y (nx19443), .A0 (nx35662), .A1 (
             camera_module_cache_ram_206__7), .S0 (nx36704)) ;
    dffr camera_module_cache_reg_ram_222__7 (.Q (camera_module_cache_ram_222__7)
         , .QB (\$dummy [2059]), .D (nx19433), .CLK (clk), .R (rst)) ;
    mux21_ni ix19434 (.Y (nx19433), .A0 (nx35662), .A1 (
             camera_module_cache_ram_222__7), .S0 (nx36708)) ;
    aoi22 ix33307 (.Y (nx33306), .A0 (camera_module_cache_ram_238__7), .A1 (
          nx37228), .B0 (camera_module_cache_ram_254__7), .B1 (nx37230)) ;
    dffr camera_module_cache_reg_ram_238__7 (.Q (camera_module_cache_ram_238__7)
         , .QB (\$dummy [2060]), .D (nx19423), .CLK (clk), .R (rst)) ;
    mux21_ni ix19424 (.Y (nx19423), .A0 (nx35664), .A1 (
             camera_module_cache_ram_238__7), .S0 (nx36712)) ;
    dffr camera_module_cache_reg_ram_254__7 (.Q (camera_module_cache_ram_254__7)
         , .QB (\$dummy [2061]), .D (nx19413), .CLK (clk), .R (rst)) ;
    mux21_ni ix19414 (.Y (nx19413), .A0 (nx35664), .A1 (
             camera_module_cache_ram_254__7), .S0 (nx36716)) ;
    oai21 ix33315 (.Y (nx33314), .A0 (nx22900), .A1 (nx22822), .B0 (nx36730)) ;
    nand04 ix22901 (.Y (nx22900), .A0 (nx33317), .A1 (nx33325), .A2 (nx33333), .A3 (
           nx33341)) ;
    aoi22 ix33318 (.Y (nx33317), .A0 (camera_module_cache_ram_15__7), .A1 (
          nx37200), .B0 (camera_module_cache_ram_31__7), .B1 (nx37202)) ;
    dffr camera_module_cache_reg_ram_15__7 (.Q (camera_module_cache_ram_15__7), 
         .QB (\$dummy [2062]), .D (nx19403), .CLK (clk), .R (rst)) ;
    mux21_ni ix19404 (.Y (nx19403), .A0 (nx35664), .A1 (
             camera_module_cache_ram_15__7), .S0 (nx36720)) ;
    dffr camera_module_cache_reg_ram_31__7 (.Q (camera_module_cache_ram_31__7), 
         .QB (\$dummy [2063]), .D (nx19393), .CLK (clk), .R (rst)) ;
    mux21_ni ix19394 (.Y (nx19393), .A0 (nx35664), .A1 (
             camera_module_cache_ram_31__7), .S0 (nx36734)) ;
    aoi22 ix33326 (.Y (nx33325), .A0 (camera_module_cache_ram_47__7), .A1 (
          nx37204), .B0 (camera_module_cache_ram_63__7), .B1 (nx37206)) ;
    dffr camera_module_cache_reg_ram_47__7 (.Q (camera_module_cache_ram_47__7), 
         .QB (\$dummy [2064]), .D (nx19383), .CLK (clk), .R (rst)) ;
    mux21_ni ix19384 (.Y (nx19383), .A0 (nx35664), .A1 (
             camera_module_cache_ram_47__7), .S0 (nx36738)) ;
    dffr camera_module_cache_reg_ram_63__7 (.Q (camera_module_cache_ram_63__7), 
         .QB (\$dummy [2065]), .D (nx19373), .CLK (clk), .R (rst)) ;
    mux21_ni ix19374 (.Y (nx19373), .A0 (nx35664), .A1 (
             camera_module_cache_ram_63__7), .S0 (nx36742)) ;
    aoi22 ix33334 (.Y (nx33333), .A0 (camera_module_cache_ram_79__7), .A1 (
          nx37208), .B0 (camera_module_cache_ram_95__7), .B1 (nx37210)) ;
    dffr camera_module_cache_reg_ram_79__7 (.Q (camera_module_cache_ram_79__7), 
         .QB (\$dummy [2066]), .D (nx19363), .CLK (clk), .R (rst)) ;
    mux21_ni ix19364 (.Y (nx19363), .A0 (nx35664), .A1 (
             camera_module_cache_ram_79__7), .S0 (nx36746)) ;
    dffr camera_module_cache_reg_ram_95__7 (.Q (camera_module_cache_ram_95__7), 
         .QB (\$dummy [2067]), .D (nx19353), .CLK (clk), .R (rst)) ;
    mux21_ni ix19354 (.Y (nx19353), .A0 (nx35666), .A1 (
             camera_module_cache_ram_95__7), .S0 (nx36750)) ;
    aoi22 ix33342 (.Y (nx33341), .A0 (camera_module_cache_ram_127__7), .A1 (
          nx37212), .B0 (camera_module_cache_ram_111__7), .B1 (nx37214)) ;
    dffr camera_module_cache_reg_ram_127__7 (.Q (camera_module_cache_ram_127__7)
         , .QB (\$dummy [2068]), .D (nx19333), .CLK (clk), .R (rst)) ;
    mux21_ni ix19334 (.Y (nx19333), .A0 (nx35666), .A1 (
             camera_module_cache_ram_127__7), .S0 (nx36754)) ;
    dffr camera_module_cache_reg_ram_111__7 (.Q (camera_module_cache_ram_111__7)
         , .QB (\$dummy [2069]), .D (nx19343), .CLK (clk), .R (rst)) ;
    mux21_ni ix19344 (.Y (nx19343), .A0 (nx35666), .A1 (
             camera_module_cache_ram_111__7), .S0 (nx36758)) ;
    nand04 ix22823 (.Y (nx22822), .A0 (nx33350), .A1 (nx33358), .A2 (nx33366), .A3 (
           nx33374)) ;
    aoi22 ix33351 (.Y (nx33350), .A0 (camera_module_cache_ram_143__7), .A1 (
          nx37216), .B0 (camera_module_cache_ram_159__7), .B1 (nx37218)) ;
    dffr camera_module_cache_reg_ram_143__7 (.Q (camera_module_cache_ram_143__7)
         , .QB (\$dummy [2070]), .D (nx19323), .CLK (clk), .R (rst)) ;
    mux21_ni ix19324 (.Y (nx19323), .A0 (nx35666), .A1 (
             camera_module_cache_ram_143__7), .S0 (nx36762)) ;
    dffr camera_module_cache_reg_ram_159__7 (.Q (camera_module_cache_ram_159__7)
         , .QB (\$dummy [2071]), .D (nx19313), .CLK (clk), .R (rst)) ;
    mux21_ni ix19314 (.Y (nx19313), .A0 (nx35666), .A1 (
             camera_module_cache_ram_159__7), .S0 (nx36766)) ;
    aoi22 ix33359 (.Y (nx33358), .A0 (camera_module_cache_ram_191__7), .A1 (
          nx37220), .B0 (camera_module_cache_ram_175__7), .B1 (nx37222)) ;
    dffr camera_module_cache_reg_ram_191__7 (.Q (camera_module_cache_ram_191__7)
         , .QB (\$dummy [2072]), .D (nx19293), .CLK (clk), .R (rst)) ;
    mux21_ni ix19294 (.Y (nx19293), .A0 (nx35666), .A1 (
             camera_module_cache_ram_191__7), .S0 (nx36770)) ;
    dffr camera_module_cache_reg_ram_175__7 (.Q (camera_module_cache_ram_175__7)
         , .QB (\$dummy [2073]), .D (nx19303), .CLK (clk), .R (rst)) ;
    mux21_ni ix19304 (.Y (nx19303), .A0 (nx35666), .A1 (
             camera_module_cache_ram_175__7), .S0 (nx36774)) ;
    aoi22 ix33367 (.Y (nx33366), .A0 (camera_module_cache_ram_207__7), .A1 (
          nx37224), .B0 (camera_module_cache_ram_223__7), .B1 (nx37226)) ;
    dffr camera_module_cache_reg_ram_207__7 (.Q (camera_module_cache_ram_207__7)
         , .QB (\$dummy [2074]), .D (nx19283), .CLK (clk), .R (rst)) ;
    mux21_ni ix19284 (.Y (nx19283), .A0 (nx35668), .A1 (
             camera_module_cache_ram_207__7), .S0 (nx36778)) ;
    dffr camera_module_cache_reg_ram_223__7 (.Q (camera_module_cache_ram_223__7)
         , .QB (\$dummy [2075]), .D (nx19273), .CLK (clk), .R (rst)) ;
    mux21_ni ix19274 (.Y (nx19273), .A0 (nx35668), .A1 (
             camera_module_cache_ram_223__7), .S0 (nx36782)) ;
    aoi22 ix33375 (.Y (nx33374), .A0 (camera_module_cache_ram_239__7), .A1 (
          nx37228), .B0 (camera_module_cache_ram_255__7), .B1 (nx37230)) ;
    dffr camera_module_cache_reg_ram_239__7 (.Q (camera_module_cache_ram_239__7)
         , .QB (\$dummy [2076]), .D (nx19263), .CLK (clk), .R (rst)) ;
    mux21_ni ix19264 (.Y (nx19263), .A0 (nx35668), .A1 (
             camera_module_cache_ram_239__7), .S0 (nx36786)) ;
    dffr camera_module_cache_reg_ram_255__7 (.Q (camera_module_cache_ram_255__7)
         , .QB (\$dummy [2077]), .D (nx19253), .CLK (clk), .R (rst)) ;
    mux21_ni ix19254 (.Y (nx19253), .A0 (nx35668), .A1 (
             camera_module_cache_ram_255__7), .S0 (nx36790)) ;
    xnor2 ix33385 (.Y (nx33384), .A0 (nx33386), .A1 (nx33472)) ;
    aoi22 ix33387 (.Y (nx33386), .A0 (zero), .A1 (nx33388), .B0 (nx26320), .B1 (
          nx26324)) ;
    oai22 ix26321 (.Y (nx26320), .A0 (nx33391), .A1 (nx33465), .B0 (nx35680), .B1 (
          nx26248)) ;
    aoi22 ix33392 (.Y (nx33391), .A0 (zero), .A1 (nx33393), .B0 (nx26172), .B1 (
          nx26176)) ;
    oai22 ix26173 (.Y (nx26172), .A0 (nx33396), .A1 (nx33458), .B0 (nx35678), .B1 (
          nx26100)) ;
    aoi22 ix33397 (.Y (nx33396), .A0 (zero), .A1 (nx33398), .B0 (nx26024), .B1 (
          nx26028)) ;
    oai22 ix26025 (.Y (nx26024), .A0 (nx33401), .A1 (nx33451), .B0 (nx35678), .B1 (
          nx25952)) ;
    aoi22 ix33402 (.Y (nx33401), .A0 (zero), .A1 (nx33403), .B0 (nx25876), .B1 (
          nx25880)) ;
    xnor2 ix33406 (.Y (nx33405), .A0 (camera_module_algo_module_pixel_value_6), 
          .A1 (nx22699)) ;
    oai22 ix25877 (.Y (nx25876), .A0 (nx33408), .A1 (nx33444), .B0 (nx35678), .B1 (
          nx25804)) ;
    aoi22 ix33409 (.Y (nx33408), .A0 (zero), .A1 (nx33410), .B0 (nx25728), .B1 (
          nx25732)) ;
    xnor2 ix33413 (.Y (nx33412), .A0 (camera_module_algo_module_pixel_value_4), 
          .A1 (nx24945)) ;
    oai22 ix25729 (.Y (nx25728), .A0 (nx33415), .A1 (nx33437), .B0 (nx35678), .B1 (
          nx25656)) ;
    aoi22 ix33416 (.Y (nx33415), .A0 (nx25580), .A1 (nx25584), .B0 (zero), .B1 (
          nx33435)) ;
    oai22 ix25581 (.Y (nx25580), .A0 (nx35678), .A1 (nx25508), .B0 (nx33419), .B1 (
          nx33427)) ;
    aoi22 ix33420 (.Y (nx33419), .A0 (one), .A1 (nx25436), .B0 (zero), .B1 (
          nx33425)) ;
    xnor2 ix25437 (.Y (nx25436), .A0 (zero), .A1 (nx25434)) ;
    xnor2 ix25435 (.Y (nx25434), .A0 (one), .A1 (nx33423)) ;
    xnor2 ix33424 (.Y (nx33423), .A0 (camera_module_algo_module_pixel_value_0), 
          .A1 (nx27681)) ;
    xnor2 ix33428 (.Y (nx33427), .A0 (zero), .A1 (nx33429)) ;
    xnor2 ix33430 (.Y (nx33429), .A0 (nx27676), .A1 (nx28817)) ;
    xnor2 ix25585 (.Y (nx25584), .A0 (zero), .A1 (nx25582)) ;
    xnor2 ix25583 (.Y (nx25582), .A0 (nx8754), .A1 (nx33433)) ;
    xnor2 ix33434 (.Y (nx33433), .A0 (camera_module_algo_module_pixel_value_2), 
          .A1 (nx26370)) ;
    xnor2 ix33438 (.Y (nx33437), .A0 (zero), .A1 (nx33439)) ;
    xnor2 ix33440 (.Y (nx33439), .A0 (nx26363), .A1 (nx29959)) ;
    xnor2 ix25733 (.Y (nx25732), .A0 (zero), .A1 (nx25730)) ;
    xnor2 ix25731 (.Y (nx25730), .A0 (nx14302), .A1 (nx33412)) ;
    xnor2 ix33445 (.Y (nx33444), .A0 (zero), .A1 (nx33446)) ;
    xnor2 ix33447 (.Y (nx33446), .A0 (nx24939), .A1 (nx31101)) ;
    xnor2 ix25881 (.Y (nx25880), .A0 (zero), .A1 (nx25878)) ;
    xnor2 ix25879 (.Y (nx25878), .A0 (nx19850), .A1 (nx33405)) ;
    xnor2 ix33452 (.Y (nx33451), .A0 (zero), .A1 (nx33453)) ;
    xnor2 ix33454 (.Y (nx33453), .A0 (nx22693), .A1 (nx32243)) ;
    xnor2 ix26029 (.Y (nx26028), .A0 (zero), .A1 (nx26026)) ;
    xnor2 ix33459 (.Y (nx33458), .A0 (zero), .A1 (nx33460)) ;
    xnor2 ix26177 (.Y (nx26176), .A0 (zero), .A1 (nx26174)) ;
    xnor2 ix33466 (.Y (nx33465), .A0 (zero), .A1 (nx33467)) ;
    xnor2 ix26325 (.Y (nx26324), .A0 (zero), .A1 (nx26322)) ;
    xnor2 ix33473 (.Y (nx33472), .A0 (zero), .A1 (nx33474)) ;
    dff camera_module_algo_module_curr_cont_reg_reg_q_13 (.Q (
        camera_module_algo_module_current_cont_value_13), .QB (nx33763), .D (
        nx22203), .CLK (clk)) ;
    dff camera_module_algo_module_Addout_reg_reg_q_13 (.Q (
        camera_module_algo_module_Addout_value_13), .QB (\$dummy [2078]), .D (
        nx22193), .CLK (clk)) ;
    xnor2 ix26359 (.Y (nx26358), .A0 (nx26356), .A1 (nx33760)) ;
    oai22 ix26357 (.Y (nx26356), .A0 (nx33485), .A1 (nx33739), .B0 (nx33753), .B1 (
          nx33750)) ;
    aoi22 ix33486 (.Y (nx33485), .A0 (camera_module_algo_module_diff_value_11), 
          .A1 (camera_module_algo_module_current_cont_value_11), .B0 (nx26208), 
          .B1 (nx929)) ;
    dff camera_module_algo_module_diff_reg_reg_q_11 (.Q (
        camera_module_algo_module_diff_value_11), .QB (nx33489), .D (nx22153), .CLK (
        clk)) ;
    aoi21 ix33492 (.Y (nx33491), .A0 (zero), .A1 (nx34122), .B0 (nx26264)) ;
    nor03_2x ix26265 (.Y (nx26264), .A0 (nx34122), .A1 (nx35700), .A2 (nx33494)
             ) ;
    xnor2 ix33495 (.Y (nx33494), .A0 (nx33391), .A1 (nx33465)) ;
    dff camera_module_algo_module_curr_cont_reg_reg_q_11 (.Q (
        camera_module_algo_module_current_cont_value_11), .QB (nx33737), .D (
        nx22143), .CLK (clk)) ;
    dff camera_module_algo_module_Addout_reg_reg_q_11 (.Q (
        camera_module_algo_module_Addout_value_11), .QB (\$dummy [2079]), .D (
        nx22133), .CLK (clk)) ;
    xnor2 ix26211 (.Y (nx26210), .A0 (nx26208), .A1 (nx33734)) ;
    oai22 ix26209 (.Y (nx26208), .A0 (nx33504), .A1 (nx33713), .B0 (nx33727), .B1 (
          nx33724)) ;
    aoi22 ix33505 (.Y (nx33504), .A0 (camera_module_algo_module_diff_value_9), .A1 (
          camera_module_algo_module_current_cont_value_9), .B0 (nx26060), .B1 (
          nx925)) ;
    dff camera_module_algo_module_diff_reg_reg_q_9 (.Q (
        camera_module_algo_module_diff_value_9), .QB (nx33508), .D (nx22093), .CLK (
        clk)) ;
    aoi21 ix33511 (.Y (nx33510), .A0 (zero), .A1 (nx34122), .B0 (nx26116)) ;
    nor03_2x ix26117 (.Y (nx26116), .A0 (nx34124), .A1 (nx35700), .A2 (nx33513)
             ) ;
    xnor2 ix33514 (.Y (nx33513), .A0 (nx33396), .A1 (nx33458)) ;
    dff camera_module_algo_module_curr_cont_reg_reg_q_9 (.Q (
        camera_module_algo_module_current_cont_value_9), .QB (nx33711), .D (
        nx22083), .CLK (clk)) ;
    dff camera_module_algo_module_Addout_reg_reg_q_9 (.Q (
        camera_module_algo_module_Addout_value_9), .QB (\$dummy [2080]), .D (
        nx22073), .CLK (clk)) ;
    xnor2 ix26063 (.Y (nx26062), .A0 (nx26060), .A1 (nx33708)) ;
    oai22 ix26061 (.Y (nx26060), .A0 (nx33523), .A1 (nx33690), .B0 (nx33707), .B1 (
          nx33701)) ;
    aoi22 ix33524 (.Y (nx33523), .A0 (camera_module_algo_module_diff_value_7), .A1 (
          camera_module_algo_module_current_cont_value_7), .B0 (nx25912), .B1 (
          nx921)) ;
    dff camera_module_algo_module_diff_reg_reg_q_7 (.Q (
        camera_module_algo_module_diff_value_7), .QB (\$dummy [2081]), .D (
        nx22033), .CLK (clk)) ;
    xnor2 ix33530 (.Y (nx33529), .A0 (nx33401), .A1 (nx33451)) ;
    dff camera_module_algo_module_curr_cont_reg_reg_q_7 (.Q (
        camera_module_algo_module_current_cont_value_7), .QB (nx33688), .D (
        nx22023), .CLK (clk)) ;
    dff camera_module_algo_module_Addout_reg_reg_q_7 (.Q (
        camera_module_algo_module_Addout_value_7), .QB (\$dummy [2082]), .D (
        nx22013), .CLK (clk)) ;
    xnor2 ix25915 (.Y (nx25914), .A0 (nx25912), .A1 (nx33685)) ;
    oai22 ix25913 (.Y (nx25912), .A0 (nx33540), .A1 (nx33667), .B0 (nx33684), .B1 (
          nx33678)) ;
    aoi22 ix33541 (.Y (nx33540), .A0 (camera_module_algo_module_diff_value_5), .A1 (
          camera_module_algo_module_current_cont_value_5), .B0 (nx25764), .B1 (
          nx917)) ;
    dff camera_module_algo_module_diff_reg_reg_q_5 (.Q (
        camera_module_algo_module_diff_value_5), .QB (\$dummy [2083]), .D (
        nx21973), .CLK (clk)) ;
    xnor2 ix33547 (.Y (nx33546), .A0 (nx33408), .A1 (nx33444)) ;
    dff camera_module_algo_module_curr_cont_reg_reg_q_5 (.Q (
        camera_module_algo_module_current_cont_value_5), .QB (nx33665), .D (
        nx21963), .CLK (clk)) ;
    dff camera_module_algo_module_Addout_reg_reg_q_5 (.Q (
        camera_module_algo_module_Addout_value_5), .QB (\$dummy [2084]), .D (
        nx21953), .CLK (clk)) ;
    xnor2 ix25767 (.Y (nx25766), .A0 (nx25764), .A1 (nx33662)) ;
    oai22 ix25765 (.Y (nx25764), .A0 (nx33557), .A1 (nx33644), .B0 (nx33661), .B1 (
          nx33655)) ;
    aoi22 ix33558 (.Y (nx33557), .A0 (camera_module_algo_module_diff_value_3), .A1 (
          camera_module_algo_module_current_cont_value_3), .B0 (nx25616), .B1 (
          nx913)) ;
    dff camera_module_algo_module_diff_reg_reg_q_3 (.Q (
        camera_module_algo_module_diff_value_3), .QB (\$dummy [2085]), .D (
        nx21913), .CLK (clk)) ;
    xnor2 ix33564 (.Y (nx33563), .A0 (nx33415), .A1 (nx33437)) ;
    dff camera_module_algo_module_curr_cont_reg_reg_q_3 (.Q (
        camera_module_algo_module_current_cont_value_3), .QB (nx33642), .D (
        nx21903), .CLK (clk)) ;
    dff camera_module_algo_module_Addout_reg_reg_q_3 (.Q (
        camera_module_algo_module_Addout_value_3), .QB (\$dummy [2086]), .D (
        nx21893), .CLK (clk)) ;
    xnor2 ix25619 (.Y (nx25618), .A0 (nx25616), .A1 (nx33639)) ;
    oai22 ix25617 (.Y (nx25616), .A0 (nx33574), .A1 (nx33621), .B0 (nx33638), .B1 (
          nx33632)) ;
    aoi22 ix33575 (.Y (nx33574), .A0 (camera_module_algo_module_diff_value_1), .A1 (
          camera_module_algo_module_current_cont_value_1), .B0 (nx25468), .B1 (
          nx910)) ;
    dff camera_module_algo_module_diff_reg_reg_q_1 (.Q (
        camera_module_algo_module_diff_value_1), .QB (\$dummy [2087]), .D (
        nx21853), .CLK (clk)) ;
    xnor2 ix33581 (.Y (nx33580), .A0 (nx33419), .A1 (nx33427)) ;
    dff camera_module_algo_module_curr_cont_reg_reg_q_1 (.Q (
        camera_module_algo_module_current_cont_value_1), .QB (nx33619), .D (
        nx21843), .CLK (clk)) ;
    dff camera_module_algo_module_Addout_reg_reg_q_1 (.Q (
        camera_module_algo_module_Addout_value_1), .QB (\$dummy [2088]), .D (
        nx21833), .CLK (clk)) ;
    xnor2 ix25471 (.Y (nx25470), .A0 (nx25468), .A1 (nx33616)) ;
    oai22 ix25469 (.Y (nx25468), .A0 (nx35680), .A1 (nx33591), .B0 (nx33615), .B1 (
          nx33609)) ;
    dff camera_module_algo_module_curr_cont_reg_reg_q_0 (.Q (
        camera_module_algo_module_current_cont_value_0), .QB (nx33609), .D (
        nx1243), .CLK (clk)) ;
    dff camera_module_algo_module_Addout_reg_reg_q_0 (.Q (
        camera_module_algo_module_Addout_value_0), .QB (\$dummy [2089]), .D (
        nx1233), .CLK (clk)) ;
    xnor2 ix657 (.Y (nx656), .A0 (zero), .A1 (nx33591)) ;
    dff camera_module_algo_module_modCU_reg_current_state_12 (.Q (
        camera_module_algo_module_modCU_current_state_12), .QB (nx33608), .D (
        nx941), .CLK (clk)) ;
    nor03_2x ix942 (.Y (nx941), .A0 (rst), .A1 (nx22979), .A2 (nx35696)) ;
    dff camera_module_algo_module_diff_reg_reg_q_0 (.Q (
        camera_module_algo_module_diff_value_0), .QB (nx33615), .D (nx21823), .CLK (
        clk)) ;
    xor2 ix25439 (.Y (nx25438), .A0 (one), .A1 (nx25436)) ;
    dff camera_module_algo_module_curr_cont_reg_reg_q_2 (.Q (
        camera_module_algo_module_current_cont_value_2), .QB (nx33632), .D (
        nx21873), .CLK (clk)) ;
    dff camera_module_algo_module_Addout_reg_reg_q_2 (.Q (
        camera_module_algo_module_Addout_value_2), .QB (\$dummy [2090]), .D (
        nx21863), .CLK (clk)) ;
    xnor2 ix33630 (.Y (nx33629), .A0 (nx33574), .A1 (nx33621)) ;
    dff camera_module_algo_module_diff_reg_reg_q_2 (.Q (
        camera_module_algo_module_diff_value_2), .QB (nx33638), .D (nx21883), .CLK (
        clk)) ;
    xor2 ix25587 (.Y (nx25586), .A0 (nx25580), .A1 (nx25584)) ;
    dff camera_module_algo_module_curr_cont_reg_reg_q_4 (.Q (
        camera_module_algo_module_current_cont_value_4), .QB (nx33655), .D (
        nx21933), .CLK (clk)) ;
    dff camera_module_algo_module_Addout_reg_reg_q_4 (.Q (
        camera_module_algo_module_Addout_value_4), .QB (\$dummy [2091]), .D (
        nx21923), .CLK (clk)) ;
    xnor2 ix33653 (.Y (nx33652), .A0 (nx33557), .A1 (nx33644)) ;
    dff camera_module_algo_module_diff_reg_reg_q_4 (.Q (
        camera_module_algo_module_diff_value_4), .QB (nx33661), .D (nx21943), .CLK (
        clk)) ;
    xor2 ix25735 (.Y (nx25734), .A0 (nx25728), .A1 (nx25732)) ;
    dff camera_module_algo_module_curr_cont_reg_reg_q_6 (.Q (
        camera_module_algo_module_current_cont_value_6), .QB (nx33678), .D (
        nx21993), .CLK (clk)) ;
    dff camera_module_algo_module_Addout_reg_reg_q_6 (.Q (
        camera_module_algo_module_Addout_value_6), .QB (\$dummy [2092]), .D (
        nx21983), .CLK (clk)) ;
    xnor2 ix33676 (.Y (nx33675), .A0 (nx33540), .A1 (nx33667)) ;
    dff camera_module_algo_module_diff_reg_reg_q_6 (.Q (
        camera_module_algo_module_diff_value_6), .QB (nx33684), .D (nx22003), .CLK (
        clk)) ;
    xor2 ix25883 (.Y (nx25882), .A0 (nx25876), .A1 (nx25880)) ;
    dff camera_module_algo_module_curr_cont_reg_reg_q_8 (.Q (
        camera_module_algo_module_current_cont_value_8), .QB (nx33701), .D (
        nx22053), .CLK (clk)) ;
    dff camera_module_algo_module_Addout_reg_reg_q_8 (.Q (
        camera_module_algo_module_Addout_value_8), .QB (\$dummy [2093]), .D (
        nx22043), .CLK (clk)) ;
    xnor2 ix33699 (.Y (nx33698), .A0 (nx33523), .A1 (nx33690)) ;
    dff camera_module_algo_module_diff_reg_reg_q_8 (.Q (
        camera_module_algo_module_diff_value_8), .QB (nx33707), .D (nx22063), .CLK (
        clk)) ;
    xor2 ix26031 (.Y (nx26030), .A0 (nx26024), .A1 (nx26028)) ;
    dff camera_module_algo_module_curr_cont_reg_reg_q_10 (.Q (
        camera_module_algo_module_current_cont_value_10), .QB (nx33724), .D (
        nx22113), .CLK (clk)) ;
    dff camera_module_algo_module_Addout_reg_reg_q_10 (.Q (
        camera_module_algo_module_Addout_value_10), .QB (\$dummy [2094]), .D (
        nx22103), .CLK (clk)) ;
    xnor2 ix33722 (.Y (nx33721), .A0 (nx33504), .A1 (nx33713)) ;
    dff camera_module_algo_module_diff_reg_reg_q_10 (.Q (\$dummy [2095]), .QB (
        nx33727), .D (nx22123), .CLK (clk)) ;
    aoi21 ix33730 (.Y (nx33729), .A0 (zero), .A1 (nx34130), .B0 (nx26190)) ;
    nor03_2x ix26191 (.Y (nx26190), .A0 (nx34130), .A1 (nx35702), .A2 (nx33732)
             ) ;
    xnor2 ix33733 (.Y (nx33732), .A0 (nx26172), .A1 (nx26176)) ;
    dff camera_module_algo_module_curr_cont_reg_reg_q_12 (.Q (
        camera_module_algo_module_current_cont_value_12), .QB (nx33750), .D (
        nx22173), .CLK (clk)) ;
    dff camera_module_algo_module_Addout_reg_reg_q_12 (.Q (
        camera_module_algo_module_Addout_value_12), .QB (\$dummy [2096]), .D (
        nx22163), .CLK (clk)) ;
    xnor2 ix33748 (.Y (nx33747), .A0 (nx33485), .A1 (nx33739)) ;
    dff camera_module_algo_module_diff_reg_reg_q_12 (.Q (\$dummy [2097]), .QB (
        nx33753), .D (nx22183), .CLK (clk)) ;
    aoi21 ix33756 (.Y (nx33755), .A0 (zero), .A1 (nx34130), .B0 (nx26338)) ;
    nor03_2x ix26339 (.Y (nx26338), .A0 (nx34130), .A1 (nx35702), .A2 (nx33758)
             ) ;
    xnor2 ix33759 (.Y (nx33758), .A0 (nx26320), .A1 (nx26324)) ;
    dff camera_module_algo_module_curr_cont_reg_reg_q_14 (.Q (
        camera_module_algo_module_current_cont_value_14), .QB (nx33776), .D (
        nx22233), .CLK (clk)) ;
    dff camera_module_algo_module_Addout_reg_reg_q_14 (.Q (
        camera_module_algo_module_Addout_value_14), .QB (\$dummy [2098]), .D (
        nx22223), .CLK (clk)) ;
    xnor2 ix33774 (.Y (nx33773), .A0 (nx22645), .A1 (nx33765)) ;
    dff camera_module_algo_module_diff_reg_reg_q_14 (.Q (\$dummy [2099]), .QB (
        nx33779), .D (nx22243), .CLK (clk)) ;
    aoi21 ix33782 (.Y (nx33781), .A0 (zero), .A1 (nx34132), .B0 (nx26486)) ;
    nor03_2x ix26487 (.Y (nx26486), .A0 (nx34132), .A1 (nx35704), .A2 (nx33784)
             ) ;
    xnor2 ix33785 (.Y (nx33784), .A0 (nx26468), .A1 (nx26472)) ;
    oai22 ix26469 (.Y (nx26468), .A0 (nx33386), .A1 (nx33472), .B0 (nx35682), .B1 (
          nx26396)) ;
    xnor2 ix26473 (.Y (nx26472), .A0 (zero), .A1 (nx26470)) ;
    dff camera_module_algo_module_diff_reg_reg_q_15 (.Q (
        camera_module_algo_module_diff_value_15), .QB (nx33794), .D (nx22253), .CLK (
        clk)) ;
    aoi21 ix33797 (.Y (nx33796), .A0 (zero), .A1 (nx34132), .B0 (nx26530)) ;
    nor03_2x ix26531 (.Y (nx26530), .A0 (nx34132), .A1 (nx35704), .A2 (nx33799)
             ) ;
    xnor2 ix33800 (.Y (nx33799), .A0 (nx33801), .A1 (nx33805)) ;
    aoi22 ix33802 (.Y (nx33801), .A0 (zero), .A1 (nx33803), .B0 (nx26468), .B1 (
          nx26472)) ;
    xnor2 ix33806 (.Y (nx33805), .A0 (zero), .A1 (nx33807)) ;
    dff camera_module_algo_module_prev_cont_reg_reg_q_15 (.Q (
        camera_module_algo_module_prev_cont_value_15), .QB (\$dummy [2100]), .D (
        nx22283), .CLK (clk)) ;
    aoi22 ix33817 (.Y (nx33816), .A0 (
          camera_module_algo_module_current_cont_value_14), .A1 (nx33818), .B0 (
          nx26604), .B1 (nx26940)) ;
    dff camera_module_algo_module_prev_cont_reg_reg_q_14 (.Q (
        camera_module_algo_module_prev_cont_value_14), .QB (nx33818), .D (
        nx22293), .CLK (clk)) ;
    oai22 ix26941 (.Y (nx26940), .A0 (nx33825), .A1 (nx33832), .B0 (nx33763), .B1 (
          camera_module_algo_module_prev_cont_value_13)) ;
    dff camera_module_algo_module_prev_cont_reg_reg_q_13 (.Q (
        camera_module_algo_module_prev_cont_value_13), .QB (\$dummy [2101]), .D (
        nx22303), .CLK (clk)) ;
    aoi22 ix33833 (.Y (nx33832), .A0 (
          camera_module_algo_module_current_cont_value_12), .A1 (nx33834), .B0 (
          nx26636), .B1 (nx26924)) ;
    dff camera_module_algo_module_prev_cont_reg_reg_q_12 (.Q (
        camera_module_algo_module_prev_cont_value_12), .QB (nx33834), .D (
        nx22313), .CLK (clk)) ;
    oai22 ix26925 (.Y (nx26924), .A0 (nx33841), .A1 (nx33848), .B0 (nx33737), .B1 (
          camera_module_algo_module_prev_cont_value_11)) ;
    dff camera_module_algo_module_prev_cont_reg_reg_q_11 (.Q (
        camera_module_algo_module_prev_cont_value_11), .QB (\$dummy [2102]), .D (
        nx22323), .CLK (clk)) ;
    aoi22 ix33849 (.Y (nx33848), .A0 (
          camera_module_algo_module_current_cont_value_10), .A1 (nx33850), .B0 (
          nx26668), .B1 (nx26908)) ;
    dff camera_module_algo_module_prev_cont_reg_reg_q_10 (.Q (
        camera_module_algo_module_prev_cont_value_10), .QB (nx33850), .D (
        nx22333), .CLK (clk)) ;
    oai22 ix26909 (.Y (nx26908), .A0 (nx33857), .A1 (nx33864), .B0 (nx33711), .B1 (
          camera_module_algo_module_prev_cont_value_9)) ;
    dff camera_module_algo_module_prev_cont_reg_reg_q_9 (.Q (
        camera_module_algo_module_prev_cont_value_9), .QB (\$dummy [2103]), .D (
        nx22343), .CLK (clk)) ;
    aoi22 ix33865 (.Y (nx33864), .A0 (
          camera_module_algo_module_current_cont_value_8), .A1 (nx33866), .B0 (
          nx26700), .B1 (nx26892)) ;
    dff camera_module_algo_module_prev_cont_reg_reg_q_8 (.Q (
        camera_module_algo_module_prev_cont_value_8), .QB (nx33866), .D (nx22353
        ), .CLK (clk)) ;
    oai22 ix26893 (.Y (nx26892), .A0 (nx33873), .A1 (nx33880), .B0 (nx33688), .B1 (
          camera_module_algo_module_prev_cont_value_7)) ;
    dff camera_module_algo_module_prev_cont_reg_reg_q_7 (.Q (
        camera_module_algo_module_prev_cont_value_7), .QB (\$dummy [2104]), .D (
        nx22363), .CLK (clk)) ;
    aoi22 ix33881 (.Y (nx33880), .A0 (
          camera_module_algo_module_current_cont_value_6), .A1 (nx33882), .B0 (
          nx26732), .B1 (nx26876)) ;
    dff camera_module_algo_module_prev_cont_reg_reg_q_6 (.Q (
        camera_module_algo_module_prev_cont_value_6), .QB (nx33882), .D (nx22373
        ), .CLK (clk)) ;
    oai22 ix26877 (.Y (nx26876), .A0 (nx33889), .A1 (nx33896), .B0 (nx33665), .B1 (
          camera_module_algo_module_prev_cont_value_5)) ;
    dff camera_module_algo_module_prev_cont_reg_reg_q_5 (.Q (
        camera_module_algo_module_prev_cont_value_5), .QB (\$dummy [2105]), .D (
        nx22383), .CLK (clk)) ;
    aoi22 ix33897 (.Y (nx33896), .A0 (
          camera_module_algo_module_current_cont_value_4), .A1 (nx33898), .B0 (
          nx26764), .B1 (nx26860)) ;
    dff camera_module_algo_module_prev_cont_reg_reg_q_4 (.Q (
        camera_module_algo_module_prev_cont_value_4), .QB (nx33898), .D (nx22393
        ), .CLK (clk)) ;
    oai22 ix26861 (.Y (nx26860), .A0 (nx33905), .A1 (nx33912), .B0 (nx33642), .B1 (
          camera_module_algo_module_prev_cont_value_3)) ;
    dff camera_module_algo_module_prev_cont_reg_reg_q_3 (.Q (
        camera_module_algo_module_prev_cont_value_3), .QB (\$dummy [2106]), .D (
        nx22403), .CLK (clk)) ;
    aoi22 ix33913 (.Y (nx33912), .A0 (
          camera_module_algo_module_current_cont_value_2), .A1 (nx33914), .B0 (
          nx26796), .B1 (nx26844)) ;
    dff camera_module_algo_module_prev_cont_reg_reg_q_2 (.Q (
        camera_module_algo_module_prev_cont_value_2), .QB (nx33914), .D (nx22413
        ), .CLK (clk)) ;
    oai22 ix26845 (.Y (nx26844), .A0 (nx33921), .A1 (nx33928), .B0 (nx33619), .B1 (
          camera_module_algo_module_prev_cont_value_1)) ;
    dff camera_module_algo_module_prev_cont_reg_reg_q_1 (.Q (
        camera_module_algo_module_prev_cont_value_1), .QB (\$dummy [2107]), .D (
        nx22423), .CLK (clk)) ;
    aoi22 ix33929 (.Y (nx33928), .A0 (
          camera_module_algo_module_current_cont_value_0), .A1 (nx33930), .B0 (
          one), .B1 (nx26828)) ;
    dff camera_module_algo_module_prev_cont_reg_reg_q_0 (.Q (
        camera_module_algo_module_prev_cont_value_0), .QB (nx33930), .D (nx22433
        ), .CLK (clk)) ;
    xnor2 ix27039 (.Y (nx27038), .A0 (
          camera_module_algo_module_current_cont_value_16), .A1 (
          camera_module_algo_module_prev_cont_value_16)) ;
    dff camera_module_algo_module_curr_cont_reg_reg_q_16 (.Q (
        camera_module_algo_module_current_cont_value_16), .QB (\$dummy [2108]), 
        .D (nx22463), .CLK (clk)) ;
    dff camera_module_algo_module_Addout_reg_reg_q_16 (.Q (
        camera_module_algo_module_Addout_value_16), .QB (\$dummy [2109]), .D (
        nx22453), .CLK (clk)) ;
    xnor2 ix33944 (.Y (nx33943), .A0 (nx33945), .A1 (nx33948)) ;
    aoi22 ix33946 (.Y (nx33945), .A0 (camera_module_algo_module_diff_value_15), 
          .A1 (camera_module_algo_module_current_cont_value_15), .B0 (nx26504), 
          .B1 (nx26542)) ;
    xnor2 ix33949 (.Y (nx33948), .A0 (
          camera_module_algo_module_current_cont_value_16), .A1 (
          camera_module_algo_module_diff_value_16)) ;
    dff camera_module_algo_module_diff_reg_reg_q_16 (.Q (
        camera_module_algo_module_diff_value_16), .QB (\$dummy [2110]), .D (
        nx22443), .CLK (clk)) ;
    oai21 ix26985 (.Y (nx26984), .A0 (nx35682), .A1 (nx35686), .B0 (nx33953)) ;
    nand03 ix33954 (.Y (nx33953), .A0 (nx26974), .A1 (nx35686), .A2 (nx37090)) ;
    xnor2 ix26975 (.Y (nx26974), .A0 (nx26970), .A1 (nx33958)) ;
    oai22 ix26971 (.Y (nx26970), .A0 (nx33801), .A1 (nx33805), .B0 (nx35682), .B1 (
          nx26514)) ;
    dff camera_module_algo_module_prev_cont_reg_reg_q_16 (.Q (
        camera_module_algo_module_prev_cont_value_16), .QB (\$dummy [2111]), .D (
        nx22473), .CLK (clk)) ;
    nand04 ix27133 (.Y (nx27132), .A0 (nx34003), .A1 (nx34005), .A2 (nx37118), .A3 (
           nx34010)) ;
    nand03 ix34006 (.Y (nx34005), .A0 (motor_move), .A1 (motor_done), .A2 (
           nx35694)) ;
    nor04 ix34011 (.Y (nx34010), .A0 (nx27122), .A1 (done), .A2 (rst), .A3 (
          nx883)) ;
    aoi21 ix27123 (.Y (nx27122), .A0 (nx22844), .A1 (nx35694), .B0 (nx22611)) ;
    dff camera_module_algo_module_modCU_reg_current_state_17 (.Q (done), .QB (
        \$dummy [2112]), .D (nx22533), .CLK (clk)) ;
    ao32 ix22534 (.Y (nx22533), .A0 (
         camera_module_algo_module_modCU_current_state_14), .A1 (nx35694), .A2 (
         camera_module_algo_module_failure_count_value_0), .B0 (done), .B1 (
         nx35696)) ;
    nor02_2x ix27121 (.Y (nx883), .A0 (rst), .A1 (nx22613)) ;
    nor03_2x ix34019 (.Y (nx34018), .A0 (nx686), .A1 (nx37082), .A2 (
             camera_module_algo_module_modCU_current_state_12)) ;
    nor02_2x ix34028 (.Y (nx34027), .A0 (done), .A1 (rst)) ;
    nand02 ix27157 (.Y (nx27156), .A0 (nx22627), .A1 (nx35686)) ;
    inv01 ix26543 (.Y (nx26542), .A (nx33790)) ;
    inv01 ix26515 (.Y (nx26514), .A (nx33807)) ;
    inv01 ix33804 (.Y (nx33803), .A (nx26470)) ;
    inv01 ix26397 (.Y (nx26396), .A (nx33474)) ;
    inv01 ix26425 (.Y (nx933), .A (nx33760)) ;
    inv01 ix33389 (.Y (nx33388), .A (nx26322)) ;
    inv01 ix26249 (.Y (nx26248), .A (nx33467)) ;
    inv01 ix26277 (.Y (nx929), .A (nx33734)) ;
    inv01 ix33394 (.Y (nx33393), .A (nx26174)) ;
    inv01 ix26101 (.Y (nx26100), .A (nx33460)) ;
    inv01 ix26129 (.Y (nx925), .A (nx33708)) ;
    inv01 ix33399 (.Y (nx33398), .A (nx26026)) ;
    inv01 ix25953 (.Y (nx25952), .A (nx33453)) ;
    inv01 ix25981 (.Y (nx921), .A (nx33685)) ;
    inv01 ix33404 (.Y (nx33403), .A (nx25878)) ;
    inv01 ix25805 (.Y (nx25804), .A (nx33446)) ;
    inv01 ix25833 (.Y (nx917), .A (nx33662)) ;
    inv01 ix33411 (.Y (nx33410), .A (nx25730)) ;
    inv01 ix25657 (.Y (nx25656), .A (nx33439)) ;
    inv01 ix25685 (.Y (nx913), .A (nx33639)) ;
    inv01 ix33436 (.Y (nx33435), .A (nx25582)) ;
    inv01 ix25509 (.Y (nx25508), .A (nx33429)) ;
    inv01 ix25537 (.Y (nx910), .A (nx33616)) ;
    inv01 ix33426 (.Y (nx33425), .A (nx25434)) ;
    inv01 ix25375 (.Y (nx25374), .A (nx32248)) ;
    inv01 ix22617 (.Y (nx22616), .A (nx33405)) ;
    inv01 ix19827 (.Y (nx19826), .A (nx31106)) ;
    inv01 ix17069 (.Y (nx17068), .A (nx33412)) ;
    inv01 ix14279 (.Y (nx14278), .A (nx29964)) ;
    inv01 ix11521 (.Y (nx11520), .A (nx33433)) ;
    inv01 ix8731 (.Y (nx8730), .A (nx28822)) ;
    inv01 ix5973 (.Y (nx5972), .A (nx33423)) ;
    inv01 ix23158 (.Y (nx23157), .A (nx986)) ;
    inv01 ix935 (.Y (nx934), .A (nx23079)) ;
    inv01 ix23530 (.Y (nx23529), .A (nx842)) ;
    inv01 ix705 (.Y (nx704), .A (nx22679)) ;
    inv01 ix585 (.Y (nx908), .A (nx23033)) ;
    inv01 ix537 (.Y (nx905), .A (nx23006)) ;
    inv01 ix479 (.Y (nx903), .A (nx22951)) ;
    inv01 ix409 (.Y (nx408), .A (nx22579)) ;
    inv01 ix405 (.Y (nx404), .A (nx22953)) ;
    inv01 ix235 (.Y (nx897), .A (nx22827)) ;
    inv01 ix129 (.Y (nx128), .A (nx22849)) ;
    inv01 ix97 (.Y (nx889), .A (nx22811)) ;
    inv02 ix34035 (.Y (nx34036), .A (nx35698)) ;
    inv02 ix34037 (.Y (nx34038), .A (nx35698)) ;
    inv02 ix34039 (.Y (nx34040), .A (nx37172)) ;
    inv02 ix34041 (.Y (nx34042), .A (nx37172)) ;
    inv02 ix34065 (.Y (nx34066), .A (nx37124)) ;
    inv02 ix34067 (.Y (nx34068), .A (nx37124)) ;
    inv02 ix34069 (.Y (nx34070), .A (nx37124)) ;
    inv02 ix34071 (.Y (nx34072), .A (nx22719)) ;
    inv02 ix34073 (.Y (nx34074), .A (nx22719)) ;
    inv02 ix34075 (.Y (nx34076), .A (nx22719)) ;
    inv02 ix34079 (.Y (nx34080), .A (nx37156)) ;
    inv02 ix34081 (.Y (nx34082), .A (nx37156)) ;
    inv02 ix34083 (.Y (nx34084), .A (nx37156)) ;
    inv02 ix34085 (.Y (nx34086), .A (nx37156)) ;
    inv02 ix34089 (.Y (nx34090), .A (nx37164)) ;
    inv02 ix34091 (.Y (nx34092), .A (nx37164)) ;
    inv02 ix34093 (.Y (nx34094), .A (nx37164)) ;
    inv02 ix34095 (.Y (nx34096), .A (nx37164)) ;
    inv02 ix34097 (.Y (nx34098), .A (nx22757)) ;
    inv02 ix34099 (.Y (nx34100), .A (nx37096)) ;
    inv02 ix34101 (.Y (nx34102), .A (nx37096)) ;
    inv02 ix34103 (.Y (nx34104), .A (nx37096)) ;
    inv02 ix34105 (.Y (nx34106), .A (nx37096)) ;
    inv02 ix34107 (.Y (nx34108), .A (nx37096)) ;
    inv02 ix34109 (.Y (nx34110), .A (nx37096)) ;
    inv02 ix34111 (.Y (nx34112), .A (nx22771)) ;
    inv02 ix34117 (.Y (nx34118), .A (nx37136)) ;
    inv02 ix34119 (.Y (nx34120), .A (nx37136)) ;
    inv02 ix34121 (.Y (nx34122), .A (nx37136)) ;
    inv02 ix34123 (.Y (nx34124), .A (nx37136)) ;
    inv02 ix34129 (.Y (nx34130), .A (nx37136)) ;
    inv02 ix34131 (.Y (nx34132), .A (nx37146)) ;
    inv02 ix34137 (.Y (nx34138), .A (nx37146)) ;
    inv04 ix34139 (.Y (nx34140), .A (nx37196)) ;
    inv04 ix34141 (.Y (nx34142), .A (nx35784)) ;
    inv02 ix34163 (.Y (nx34164), .A (nx36804)) ;
    inv02 ix34165 (.Y (nx34166), .A (nx36804)) ;
    inv02 ix34167 (.Y (nx34168), .A (nx36804)) ;
    inv02 ix34169 (.Y (nx34170), .A (nx36804)) ;
    inv02 ix34171 (.Y (nx34172), .A (nx36804)) ;
    inv02 ix34173 (.Y (nx34174), .A (nx36804)) ;
    inv02 ix34175 (.Y (nx34176), .A (nx36804)) ;
    inv02 ix34177 (.Y (nx34178), .A (nx36806)) ;
    inv02 ix34179 (.Y (nx34180), .A (nx36806)) ;
    inv02 ix34181 (.Y (nx34182), .A (nx36806)) ;
    inv02 ix34183 (.Y (nx34184), .A (nx36806)) ;
    inv02 ix34185 (.Y (nx34186), .A (nx36806)) ;
    inv02 ix34187 (.Y (nx34188), .A (nx36806)) ;
    inv02 ix34189 (.Y (nx34190), .A (nx36806)) ;
    inv02 ix34191 (.Y (nx34192), .A (nx36808)) ;
    inv02 ix34193 (.Y (nx34194), .A (nx36808)) ;
    inv02 ix34195 (.Y (nx34196), .A (nx36808)) ;
    inv02 ix34197 (.Y (nx34198), .A (nx36808)) ;
    inv02 ix34199 (.Y (nx34200), .A (nx36808)) ;
    inv02 ix34201 (.Y (nx34202), .A (nx36808)) ;
    inv02 ix34203 (.Y (nx34204), .A (nx36808)) ;
    inv02 ix34205 (.Y (nx34206), .A (nx36810)) ;
    inv02 ix34207 (.Y (nx34208), .A (nx36810)) ;
    inv02 ix34209 (.Y (nx34210), .A (nx36810)) ;
    inv02 ix34211 (.Y (nx34212), .A (nx36810)) ;
    inv02 ix34213 (.Y (nx34214), .A (nx36810)) ;
    inv02 ix34215 (.Y (nx34216), .A (nx36810)) ;
    inv02 ix34217 (.Y (nx34218), .A (nx36810)) ;
    inv02 ix34219 (.Y (nx34220), .A (nx36812)) ;
    inv02 ix34221 (.Y (nx34222), .A (nx36812)) ;
    inv02 ix34223 (.Y (nx34224), .A (nx36812)) ;
    inv02 ix34225 (.Y (nx34226), .A (nx36812)) ;
    inv02 ix34227 (.Y (nx34228), .A (nx36812)) ;
    inv02 ix34229 (.Y (nx34230), .A (nx36812)) ;
    inv02 ix34231 (.Y (nx34232), .A (nx36812)) ;
    inv02 ix34233 (.Y (nx34234), .A (nx36814)) ;
    inv02 ix34235 (.Y (nx34236), .A (nx36814)) ;
    buf02 ix34303 (.Y (nx34304), .A (nx2424)) ;
    buf02 ix34305 (.Y (nx34306), .A (nx2424)) ;
    buf02 ix34307 (.Y (nx34308), .A (nx2440)) ;
    buf02 ix34309 (.Y (nx34310), .A (nx2440)) ;
    buf02 ix34311 (.Y (nx34312), .A (nx2458)) ;
    buf02 ix34313 (.Y (nx34314), .A (nx2458)) ;
    buf02 ix34315 (.Y (nx34316), .A (nx2474)) ;
    buf02 ix34317 (.Y (nx34318), .A (nx2474)) ;
    buf02 ix34319 (.Y (nx34320), .A (nx2494)) ;
    buf02 ix34321 (.Y (nx34322), .A (nx2494)) ;
    buf02 ix34323 (.Y (nx34324), .A (nx2510)) ;
    buf02 ix34325 (.Y (nx34326), .A (nx2510)) ;
    buf02 ix34327 (.Y (nx34328), .A (nx2528)) ;
    buf02 ix34329 (.Y (nx34330), .A (nx2528)) ;
    buf02 ix34331 (.Y (nx34332), .A (nx2544)) ;
    buf02 ix34333 (.Y (nx34334), .A (nx2544)) ;
    buf02 ix34335 (.Y (nx34336), .A (nx2566)) ;
    buf02 ix34337 (.Y (nx34338), .A (nx2566)) ;
    buf02 ix34339 (.Y (nx34340), .A (nx2582)) ;
    buf02 ix34341 (.Y (nx34342), .A (nx2582)) ;
    buf02 ix34343 (.Y (nx34344), .A (nx2600)) ;
    buf02 ix34345 (.Y (nx34346), .A (nx2600)) ;
    buf02 ix34347 (.Y (nx34348), .A (nx2616)) ;
    buf02 ix34349 (.Y (nx34350), .A (nx2616)) ;
    buf02 ix34351 (.Y (nx34352), .A (nx2636)) ;
    buf02 ix34353 (.Y (nx34354), .A (nx2636)) ;
    buf02 ix34355 (.Y (nx34356), .A (nx2652)) ;
    buf02 ix34357 (.Y (nx34358), .A (nx2652)) ;
    buf02 ix34359 (.Y (nx34360), .A (nx2670)) ;
    buf02 ix34361 (.Y (nx34362), .A (nx2670)) ;
    buf02 ix34363 (.Y (nx34364), .A (nx2686)) ;
    buf02 ix34365 (.Y (nx34366), .A (nx2686)) ;
    buf02 ix34373 (.Y (nx34374), .A (nx2716)) ;
    buf02 ix34375 (.Y (nx34376), .A (nx2716)) ;
    buf02 ix34377 (.Y (nx34378), .A (nx2732)) ;
    buf02 ix34379 (.Y (nx34380), .A (nx2732)) ;
    buf02 ix34381 (.Y (nx34382), .A (nx2750)) ;
    buf02 ix34383 (.Y (nx34384), .A (nx2750)) ;
    buf02 ix34385 (.Y (nx34386), .A (nx2766)) ;
    buf02 ix34387 (.Y (nx34388), .A (nx2766)) ;
    buf02 ix34389 (.Y (nx34390), .A (nx2786)) ;
    buf02 ix34391 (.Y (nx34392), .A (nx2786)) ;
    buf02 ix34393 (.Y (nx34394), .A (nx2802)) ;
    buf02 ix34395 (.Y (nx34396), .A (nx2802)) ;
    buf02 ix34397 (.Y (nx34398), .A (nx2820)) ;
    buf02 ix34399 (.Y (nx34400), .A (nx2820)) ;
    buf02 ix34401 (.Y (nx34402), .A (nx2836)) ;
    buf02 ix34403 (.Y (nx34404), .A (nx2836)) ;
    buf02 ix34405 (.Y (nx34406), .A (nx2858)) ;
    buf02 ix34407 (.Y (nx34408), .A (nx2858)) ;
    buf02 ix34409 (.Y (nx34410), .A (nx2874)) ;
    buf02 ix34411 (.Y (nx34412), .A (nx2874)) ;
    buf02 ix34413 (.Y (nx34414), .A (nx2892)) ;
    buf02 ix34415 (.Y (nx34416), .A (nx2892)) ;
    buf02 ix34417 (.Y (nx34418), .A (nx2908)) ;
    buf02 ix34419 (.Y (nx34420), .A (nx2908)) ;
    buf02 ix34421 (.Y (nx34422), .A (nx2928)) ;
    buf02 ix34423 (.Y (nx34424), .A (nx2928)) ;
    buf02 ix34425 (.Y (nx34426), .A (nx2944)) ;
    buf02 ix34427 (.Y (nx34428), .A (nx2944)) ;
    buf02 ix34429 (.Y (nx34430), .A (nx2962)) ;
    buf02 ix34431 (.Y (nx34432), .A (nx2962)) ;
    buf02 ix34433 (.Y (nx34434), .A (nx2978)) ;
    buf02 ix34435 (.Y (nx34436), .A (nx2978)) ;
    buf02 ix34443 (.Y (nx34444), .A (nx3010)) ;
    buf02 ix34445 (.Y (nx34446), .A (nx3010)) ;
    buf02 ix34447 (.Y (nx34448), .A (nx3026)) ;
    buf02 ix34449 (.Y (nx34450), .A (nx3026)) ;
    buf02 ix34451 (.Y (nx34452), .A (nx3044)) ;
    buf02 ix34453 (.Y (nx34454), .A (nx3044)) ;
    buf02 ix34455 (.Y (nx34456), .A (nx3060)) ;
    buf02 ix34457 (.Y (nx34458), .A (nx3060)) ;
    buf02 ix34459 (.Y (nx34460), .A (nx3080)) ;
    buf02 ix34461 (.Y (nx34462), .A (nx3080)) ;
    buf02 ix34463 (.Y (nx34464), .A (nx3096)) ;
    buf02 ix34465 (.Y (nx34466), .A (nx3096)) ;
    buf02 ix34467 (.Y (nx34468), .A (nx3114)) ;
    buf02 ix34469 (.Y (nx34470), .A (nx3114)) ;
    buf02 ix34471 (.Y (nx34472), .A (nx3130)) ;
    buf02 ix34473 (.Y (nx34474), .A (nx3130)) ;
    buf02 ix34475 (.Y (nx34476), .A (nx3152)) ;
    buf02 ix34477 (.Y (nx34478), .A (nx3152)) ;
    buf02 ix34479 (.Y (nx34480), .A (nx3168)) ;
    buf02 ix34481 (.Y (nx34482), .A (nx3168)) ;
    buf02 ix34483 (.Y (nx34484), .A (nx3186)) ;
    buf02 ix34485 (.Y (nx34486), .A (nx3186)) ;
    buf02 ix34487 (.Y (nx34488), .A (nx3202)) ;
    buf02 ix34489 (.Y (nx34490), .A (nx3202)) ;
    buf02 ix34491 (.Y (nx34492), .A (nx3222)) ;
    buf02 ix34493 (.Y (nx34494), .A (nx3222)) ;
    buf02 ix34495 (.Y (nx34496), .A (nx3238)) ;
    buf02 ix34497 (.Y (nx34498), .A (nx3238)) ;
    buf02 ix34499 (.Y (nx34500), .A (nx3256)) ;
    buf02 ix34501 (.Y (nx34502), .A (nx3256)) ;
    buf02 ix34503 (.Y (nx34504), .A (nx3272)) ;
    buf02 ix34505 (.Y (nx34506), .A (nx3272)) ;
    buf02 ix34513 (.Y (nx34514), .A (nx3302)) ;
    buf02 ix34515 (.Y (nx34516), .A (nx3302)) ;
    buf02 ix34517 (.Y (nx34518), .A (nx3318)) ;
    buf02 ix34519 (.Y (nx34520), .A (nx3318)) ;
    buf02 ix34521 (.Y (nx34522), .A (nx3336)) ;
    buf02 ix34523 (.Y (nx34524), .A (nx3336)) ;
    buf02 ix34525 (.Y (nx34526), .A (nx3352)) ;
    buf02 ix34527 (.Y (nx34528), .A (nx3352)) ;
    buf02 ix34529 (.Y (nx34530), .A (nx3372)) ;
    buf02 ix34531 (.Y (nx34532), .A (nx3372)) ;
    buf02 ix34533 (.Y (nx34534), .A (nx3388)) ;
    buf02 ix34535 (.Y (nx34536), .A (nx3388)) ;
    buf02 ix34537 (.Y (nx34538), .A (nx3406)) ;
    buf02 ix34539 (.Y (nx34540), .A (nx3406)) ;
    buf02 ix34541 (.Y (nx34542), .A (nx3422)) ;
    buf02 ix34543 (.Y (nx34544), .A (nx3422)) ;
    buf02 ix34545 (.Y (nx34546), .A (nx3444)) ;
    buf02 ix34547 (.Y (nx34548), .A (nx3444)) ;
    buf02 ix34549 (.Y (nx34550), .A (nx3460)) ;
    buf02 ix34551 (.Y (nx34552), .A (nx3460)) ;
    buf02 ix34553 (.Y (nx34554), .A (nx3478)) ;
    buf02 ix34555 (.Y (nx34556), .A (nx3478)) ;
    buf02 ix34557 (.Y (nx34558), .A (nx3494)) ;
    buf02 ix34559 (.Y (nx34560), .A (nx3494)) ;
    buf02 ix34561 (.Y (nx34562), .A (nx3514)) ;
    buf02 ix34563 (.Y (nx34564), .A (nx3514)) ;
    buf02 ix34565 (.Y (nx34566), .A (nx3530)) ;
    buf02 ix34567 (.Y (nx34568), .A (nx3530)) ;
    buf02 ix34569 (.Y (nx34570), .A (nx3548)) ;
    buf02 ix34571 (.Y (nx34572), .A (nx3548)) ;
    buf02 ix34573 (.Y (nx34574), .A (nx3564)) ;
    buf02 ix34575 (.Y (nx34576), .A (nx3564)) ;
    buf02 ix34583 (.Y (nx34584), .A (nx3604)) ;
    buf02 ix34585 (.Y (nx34586), .A (nx3604)) ;
    buf02 ix34587 (.Y (nx34588), .A (nx3620)) ;
    buf02 ix34589 (.Y (nx34590), .A (nx3620)) ;
    buf02 ix34591 (.Y (nx34592), .A (nx3638)) ;
    buf02 ix34593 (.Y (nx34594), .A (nx3638)) ;
    buf02 ix34595 (.Y (nx34596), .A (nx3654)) ;
    buf02 ix34597 (.Y (nx34598), .A (nx3654)) ;
    buf02 ix34599 (.Y (nx34600), .A (nx3674)) ;
    buf02 ix34601 (.Y (nx34602), .A (nx3674)) ;
    buf02 ix34603 (.Y (nx34604), .A (nx3690)) ;
    buf02 ix34605 (.Y (nx34606), .A (nx3690)) ;
    buf02 ix34607 (.Y (nx34608), .A (nx3708)) ;
    buf02 ix34609 (.Y (nx34610), .A (nx3708)) ;
    buf02 ix34611 (.Y (nx34612), .A (nx3724)) ;
    buf02 ix34613 (.Y (nx34614), .A (nx3724)) ;
    buf02 ix34615 (.Y (nx34616), .A (nx3746)) ;
    buf02 ix34617 (.Y (nx34618), .A (nx3746)) ;
    buf02 ix34619 (.Y (nx34620), .A (nx3762)) ;
    buf02 ix34621 (.Y (nx34622), .A (nx3762)) ;
    buf02 ix34623 (.Y (nx34624), .A (nx3780)) ;
    buf02 ix34625 (.Y (nx34626), .A (nx3780)) ;
    buf02 ix34627 (.Y (nx34628), .A (nx3796)) ;
    buf02 ix34629 (.Y (nx34630), .A (nx3796)) ;
    buf02 ix34631 (.Y (nx34632), .A (nx3816)) ;
    buf02 ix34633 (.Y (nx34634), .A (nx3816)) ;
    buf02 ix34635 (.Y (nx34636), .A (nx3832)) ;
    buf02 ix34637 (.Y (nx34638), .A (nx3832)) ;
    buf02 ix34639 (.Y (nx34640), .A (nx3850)) ;
    buf02 ix34641 (.Y (nx34642), .A (nx3850)) ;
    buf02 ix34643 (.Y (nx34644), .A (nx3866)) ;
    buf02 ix34645 (.Y (nx34646), .A (nx3866)) ;
    buf02 ix34653 (.Y (nx34654), .A (nx3896)) ;
    buf02 ix34655 (.Y (nx34656), .A (nx3896)) ;
    buf02 ix34657 (.Y (nx34658), .A (nx3912)) ;
    buf02 ix34659 (.Y (nx34660), .A (nx3912)) ;
    buf02 ix34661 (.Y (nx34662), .A (nx3930)) ;
    buf02 ix34663 (.Y (nx34664), .A (nx3930)) ;
    buf02 ix34665 (.Y (nx34666), .A (nx3946)) ;
    buf02 ix34667 (.Y (nx34668), .A (nx3946)) ;
    buf02 ix34669 (.Y (nx34670), .A (nx3966)) ;
    buf02 ix34671 (.Y (nx34672), .A (nx3966)) ;
    buf02 ix34673 (.Y (nx34674), .A (nx3982)) ;
    buf02 ix34675 (.Y (nx34676), .A (nx3982)) ;
    buf02 ix34677 (.Y (nx34678), .A (nx4000)) ;
    buf02 ix34679 (.Y (nx34680), .A (nx4000)) ;
    buf02 ix34681 (.Y (nx34682), .A (nx4016)) ;
    buf02 ix34683 (.Y (nx34684), .A (nx4016)) ;
    buf02 ix34685 (.Y (nx34686), .A (nx4038)) ;
    buf02 ix34687 (.Y (nx34688), .A (nx4038)) ;
    buf02 ix34689 (.Y (nx34690), .A (nx4054)) ;
    buf02 ix34691 (.Y (nx34692), .A (nx4054)) ;
    buf02 ix34693 (.Y (nx34694), .A (nx4072)) ;
    buf02 ix34695 (.Y (nx34696), .A (nx4072)) ;
    buf02 ix34697 (.Y (nx34698), .A (nx4088)) ;
    buf02 ix34699 (.Y (nx34700), .A (nx4088)) ;
    buf02 ix34701 (.Y (nx34702), .A (nx4108)) ;
    buf02 ix34703 (.Y (nx34704), .A (nx4108)) ;
    buf02 ix34705 (.Y (nx34706), .A (nx4124)) ;
    buf02 ix34707 (.Y (nx34708), .A (nx4124)) ;
    buf02 ix34709 (.Y (nx34710), .A (nx4142)) ;
    buf02 ix34711 (.Y (nx34712), .A (nx4142)) ;
    buf02 ix34713 (.Y (nx34714), .A (nx4158)) ;
    buf02 ix34715 (.Y (nx34716), .A (nx4158)) ;
    buf02 ix34723 (.Y (nx34724), .A (nx4190)) ;
    buf02 ix34725 (.Y (nx34726), .A (nx4190)) ;
    buf02 ix34727 (.Y (nx34728), .A (nx4206)) ;
    buf02 ix34729 (.Y (nx34730), .A (nx4206)) ;
    buf02 ix34731 (.Y (nx34732), .A (nx4224)) ;
    buf02 ix34733 (.Y (nx34734), .A (nx4224)) ;
    buf02 ix34735 (.Y (nx34736), .A (nx4240)) ;
    buf02 ix34737 (.Y (nx34738), .A (nx4240)) ;
    buf02 ix34739 (.Y (nx34740), .A (nx4260)) ;
    buf02 ix34741 (.Y (nx34742), .A (nx4260)) ;
    buf02 ix34743 (.Y (nx34744), .A (nx4276)) ;
    buf02 ix34745 (.Y (nx34746), .A (nx4276)) ;
    buf02 ix34747 (.Y (nx34748), .A (nx4294)) ;
    buf02 ix34749 (.Y (nx34750), .A (nx4294)) ;
    buf02 ix34751 (.Y (nx34752), .A (nx4310)) ;
    buf02 ix34753 (.Y (nx34754), .A (nx4310)) ;
    buf02 ix34755 (.Y (nx34756), .A (nx4332)) ;
    buf02 ix34757 (.Y (nx34758), .A (nx4332)) ;
    buf02 ix34759 (.Y (nx34760), .A (nx4348)) ;
    buf02 ix34761 (.Y (nx34762), .A (nx4348)) ;
    buf02 ix34763 (.Y (nx34764), .A (nx4366)) ;
    buf02 ix34765 (.Y (nx34766), .A (nx4366)) ;
    buf02 ix34767 (.Y (nx34768), .A (nx4382)) ;
    buf02 ix34769 (.Y (nx34770), .A (nx4382)) ;
    buf02 ix34771 (.Y (nx34772), .A (nx4402)) ;
    buf02 ix34773 (.Y (nx34774), .A (nx4402)) ;
    buf02 ix34775 (.Y (nx34776), .A (nx4418)) ;
    buf02 ix34777 (.Y (nx34778), .A (nx4418)) ;
    buf02 ix34779 (.Y (nx34780), .A (nx4436)) ;
    buf02 ix34781 (.Y (nx34782), .A (nx4436)) ;
    buf02 ix34783 (.Y (nx34784), .A (nx4452)) ;
    buf02 ix34785 (.Y (nx34786), .A (nx4452)) ;
    buf02 ix34793 (.Y (nx34794), .A (nx4482)) ;
    buf02 ix34795 (.Y (nx34796), .A (nx4482)) ;
    buf02 ix34797 (.Y (nx34798), .A (nx4498)) ;
    buf02 ix34799 (.Y (nx34800), .A (nx4498)) ;
    buf02 ix34801 (.Y (nx34802), .A (nx4516)) ;
    buf02 ix34803 (.Y (nx34804), .A (nx4516)) ;
    buf02 ix34805 (.Y (nx34806), .A (nx4532)) ;
    buf02 ix34807 (.Y (nx34808), .A (nx4532)) ;
    buf02 ix34809 (.Y (nx34810), .A (nx4552)) ;
    buf02 ix34811 (.Y (nx34812), .A (nx4552)) ;
    buf02 ix34813 (.Y (nx34814), .A (nx4568)) ;
    buf02 ix34815 (.Y (nx34816), .A (nx4568)) ;
    buf02 ix34817 (.Y (nx34818), .A (nx4586)) ;
    buf02 ix34819 (.Y (nx34820), .A (nx4586)) ;
    buf02 ix34821 (.Y (nx34822), .A (nx4602)) ;
    buf02 ix34823 (.Y (nx34824), .A (nx4602)) ;
    buf02 ix34825 (.Y (nx34826), .A (nx4624)) ;
    buf02 ix34827 (.Y (nx34828), .A (nx4624)) ;
    buf02 ix34829 (.Y (nx34830), .A (nx4640)) ;
    buf02 ix34831 (.Y (nx34832), .A (nx4640)) ;
    buf02 ix34833 (.Y (nx34834), .A (nx4658)) ;
    buf02 ix34835 (.Y (nx34836), .A (nx4658)) ;
    buf02 ix34837 (.Y (nx34838), .A (nx4674)) ;
    buf02 ix34839 (.Y (nx34840), .A (nx4674)) ;
    buf02 ix34841 (.Y (nx34842), .A (nx4694)) ;
    buf02 ix34843 (.Y (nx34844), .A (nx4694)) ;
    buf02 ix34845 (.Y (nx34846), .A (nx4710)) ;
    buf02 ix34847 (.Y (nx34848), .A (nx4710)) ;
    buf02 ix34849 (.Y (nx34850), .A (nx4728)) ;
    buf02 ix34851 (.Y (nx34852), .A (nx4728)) ;
    buf02 ix34853 (.Y (nx34854), .A (nx4744)) ;
    buf02 ix34855 (.Y (nx34856), .A (nx4744)) ;
    buf02 ix34863 (.Y (nx34864), .A (nx4780)) ;
    buf02 ix34865 (.Y (nx34866), .A (nx4780)) ;
    buf02 ix34867 (.Y (nx34868), .A (nx4796)) ;
    buf02 ix34869 (.Y (nx34870), .A (nx4796)) ;
    buf02 ix34871 (.Y (nx34872), .A (nx4814)) ;
    buf02 ix34873 (.Y (nx34874), .A (nx4814)) ;
    buf02 ix34875 (.Y (nx34876), .A (nx4830)) ;
    buf02 ix34877 (.Y (nx34878), .A (nx4830)) ;
    buf02 ix34879 (.Y (nx34880), .A (nx4850)) ;
    buf02 ix34881 (.Y (nx34882), .A (nx4850)) ;
    buf02 ix34883 (.Y (nx34884), .A (nx4866)) ;
    buf02 ix34885 (.Y (nx34886), .A (nx4866)) ;
    buf02 ix34887 (.Y (nx34888), .A (nx4884)) ;
    buf02 ix34889 (.Y (nx34890), .A (nx4884)) ;
    buf02 ix34891 (.Y (nx34892), .A (nx4900)) ;
    buf02 ix34893 (.Y (nx34894), .A (nx4900)) ;
    buf02 ix34895 (.Y (nx34896), .A (nx4922)) ;
    buf02 ix34897 (.Y (nx34898), .A (nx4922)) ;
    buf02 ix34899 (.Y (nx34900), .A (nx4938)) ;
    buf02 ix34901 (.Y (nx34902), .A (nx4938)) ;
    buf02 ix34903 (.Y (nx34904), .A (nx4956)) ;
    buf02 ix34905 (.Y (nx34906), .A (nx4956)) ;
    buf02 ix34907 (.Y (nx34908), .A (nx4972)) ;
    buf02 ix34909 (.Y (nx34910), .A (nx4972)) ;
    buf02 ix34911 (.Y (nx34912), .A (nx4992)) ;
    buf02 ix34913 (.Y (nx34914), .A (nx4992)) ;
    buf02 ix34915 (.Y (nx34916), .A (nx5008)) ;
    buf02 ix34917 (.Y (nx34918), .A (nx5008)) ;
    buf02 ix34919 (.Y (nx34920), .A (nx5026)) ;
    buf02 ix34921 (.Y (nx34922), .A (nx5026)) ;
    buf02 ix34923 (.Y (nx34924), .A (nx5042)) ;
    buf02 ix34925 (.Y (nx34926), .A (nx5042)) ;
    buf02 ix34933 (.Y (nx34934), .A (nx5072)) ;
    buf02 ix34935 (.Y (nx34936), .A (nx5072)) ;
    buf02 ix34937 (.Y (nx34938), .A (nx5088)) ;
    buf02 ix34939 (.Y (nx34940), .A (nx5088)) ;
    buf02 ix34941 (.Y (nx34942), .A (nx5106)) ;
    buf02 ix34943 (.Y (nx34944), .A (nx5106)) ;
    buf02 ix34945 (.Y (nx34946), .A (nx5122)) ;
    buf02 ix34947 (.Y (nx34948), .A (nx5122)) ;
    buf02 ix34949 (.Y (nx34950), .A (nx5142)) ;
    buf02 ix34951 (.Y (nx34952), .A (nx5142)) ;
    buf02 ix34953 (.Y (nx34954), .A (nx5158)) ;
    buf02 ix34955 (.Y (nx34956), .A (nx5158)) ;
    buf02 ix34957 (.Y (nx34958), .A (nx5176)) ;
    buf02 ix34959 (.Y (nx34960), .A (nx5176)) ;
    buf02 ix34961 (.Y (nx34962), .A (nx5192)) ;
    buf02 ix34963 (.Y (nx34964), .A (nx5192)) ;
    buf02 ix34965 (.Y (nx34966), .A (nx5214)) ;
    buf02 ix34967 (.Y (nx34968), .A (nx5214)) ;
    buf02 ix34969 (.Y (nx34970), .A (nx5230)) ;
    buf02 ix34971 (.Y (nx34972), .A (nx5230)) ;
    buf02 ix34973 (.Y (nx34974), .A (nx5248)) ;
    buf02 ix34975 (.Y (nx34976), .A (nx5248)) ;
    buf02 ix34977 (.Y (nx34978), .A (nx5264)) ;
    buf02 ix34979 (.Y (nx34980), .A (nx5264)) ;
    buf02 ix34981 (.Y (nx34982), .A (nx5284)) ;
    buf02 ix34983 (.Y (nx34984), .A (nx5284)) ;
    buf02 ix34985 (.Y (nx34986), .A (nx5300)) ;
    buf02 ix34987 (.Y (nx34988), .A (nx5300)) ;
    buf02 ix34989 (.Y (nx34990), .A (nx5318)) ;
    buf02 ix34991 (.Y (nx34992), .A (nx5318)) ;
    buf02 ix34993 (.Y (nx34994), .A (nx5334)) ;
    buf02 ix34995 (.Y (nx34996), .A (nx5334)) ;
    buf02 ix35003 (.Y (nx35004), .A (nx5366)) ;
    buf02 ix35005 (.Y (nx35006), .A (nx5366)) ;
    buf02 ix35007 (.Y (nx35008), .A (nx5382)) ;
    buf02 ix35009 (.Y (nx35010), .A (nx5382)) ;
    buf02 ix35011 (.Y (nx35012), .A (nx5400)) ;
    buf02 ix35013 (.Y (nx35014), .A (nx5400)) ;
    buf02 ix35015 (.Y (nx35016), .A (nx5416)) ;
    buf02 ix35017 (.Y (nx35018), .A (nx5416)) ;
    buf02 ix35019 (.Y (nx35020), .A (nx5436)) ;
    buf02 ix35021 (.Y (nx35022), .A (nx5436)) ;
    buf02 ix35023 (.Y (nx35024), .A (nx5452)) ;
    buf02 ix35025 (.Y (nx35026), .A (nx5452)) ;
    buf02 ix35027 (.Y (nx35028), .A (nx5470)) ;
    buf02 ix35029 (.Y (nx35030), .A (nx5470)) ;
    buf02 ix35031 (.Y (nx35032), .A (nx5486)) ;
    buf02 ix35033 (.Y (nx35034), .A (nx5486)) ;
    buf02 ix35035 (.Y (nx35036), .A (nx5508)) ;
    buf02 ix35037 (.Y (nx35038), .A (nx5508)) ;
    buf02 ix35039 (.Y (nx35040), .A (nx5524)) ;
    buf02 ix35041 (.Y (nx35042), .A (nx5524)) ;
    buf02 ix35043 (.Y (nx35044), .A (nx5542)) ;
    buf02 ix35045 (.Y (nx35046), .A (nx5542)) ;
    buf02 ix35047 (.Y (nx35048), .A (nx5558)) ;
    buf02 ix35049 (.Y (nx35050), .A (nx5558)) ;
    buf02 ix35051 (.Y (nx35052), .A (nx5578)) ;
    buf02 ix35053 (.Y (nx35054), .A (nx5578)) ;
    buf02 ix35055 (.Y (nx35056), .A (nx5594)) ;
    buf02 ix35057 (.Y (nx35058), .A (nx5594)) ;
    buf02 ix35059 (.Y (nx35060), .A (nx5612)) ;
    buf02 ix35061 (.Y (nx35062), .A (nx5612)) ;
    buf02 ix35063 (.Y (nx35064), .A (nx5628)) ;
    buf02 ix35065 (.Y (nx35066), .A (nx5628)) ;
    buf02 ix35073 (.Y (nx35074), .A (nx5658)) ;
    buf02 ix35075 (.Y (nx35076), .A (nx5658)) ;
    buf02 ix35077 (.Y (nx35078), .A (nx5674)) ;
    buf02 ix35079 (.Y (nx35080), .A (nx5674)) ;
    buf02 ix35081 (.Y (nx35082), .A (nx5692)) ;
    buf02 ix35083 (.Y (nx35084), .A (nx5692)) ;
    buf02 ix35085 (.Y (nx35086), .A (nx5708)) ;
    buf02 ix35087 (.Y (nx35088), .A (nx5708)) ;
    buf02 ix35089 (.Y (nx35090), .A (nx5728)) ;
    buf02 ix35091 (.Y (nx35092), .A (nx5728)) ;
    buf02 ix35093 (.Y (nx35094), .A (nx5744)) ;
    buf02 ix35095 (.Y (nx35096), .A (nx5744)) ;
    buf02 ix35097 (.Y (nx35098), .A (nx5762)) ;
    buf02 ix35099 (.Y (nx35100), .A (nx5762)) ;
    buf02 ix35101 (.Y (nx35102), .A (nx5778)) ;
    buf02 ix35103 (.Y (nx35104), .A (nx5778)) ;
    buf02 ix35105 (.Y (nx35106), .A (nx5800)) ;
    buf02 ix35107 (.Y (nx35108), .A (nx5800)) ;
    buf02 ix35109 (.Y (nx35110), .A (nx5816)) ;
    buf02 ix35111 (.Y (nx35112), .A (nx5816)) ;
    buf02 ix35113 (.Y (nx35114), .A (nx5834)) ;
    buf02 ix35115 (.Y (nx35116), .A (nx5834)) ;
    buf02 ix35117 (.Y (nx35118), .A (nx5850)) ;
    buf02 ix35119 (.Y (nx35120), .A (nx5850)) ;
    buf02 ix35121 (.Y (nx35122), .A (nx5870)) ;
    buf02 ix35123 (.Y (nx35124), .A (nx5870)) ;
    buf02 ix35125 (.Y (nx35126), .A (nx5886)) ;
    buf02 ix35127 (.Y (nx35128), .A (nx5886)) ;
    buf02 ix35129 (.Y (nx35130), .A (nx5904)) ;
    buf02 ix35131 (.Y (nx35132), .A (nx5904)) ;
    buf02 ix35133 (.Y (nx35134), .A (nx5920)) ;
    buf02 ix35135 (.Y (nx35136), .A (nx5920)) ;
    inv02 ix35139 (.Y (nx35140), .A (nx36816)) ;
    inv02 ix35141 (.Y (nx35142), .A (nx36816)) ;
    inv02 ix35143 (.Y (nx35144), .A (nx36816)) ;
    inv02 ix35145 (.Y (nx35146), .A (nx36816)) ;
    inv02 ix35147 (.Y (nx35148), .A (nx36816)) ;
    inv02 ix35149 (.Y (nx35150), .A (nx36816)) ;
    inv02 ix35151 (.Y (nx35152), .A (nx36816)) ;
    inv02 ix35153 (.Y (nx35154), .A (nx36818)) ;
    inv02 ix35155 (.Y (nx35156), .A (nx36818)) ;
    inv02 ix35157 (.Y (nx35158), .A (nx36818)) ;
    inv02 ix35159 (.Y (nx35160), .A (nx36818)) ;
    inv02 ix35161 (.Y (nx35162), .A (nx36818)) ;
    inv02 ix35163 (.Y (nx35164), .A (nx36818)) ;
    inv02 ix35165 (.Y (nx35166), .A (nx36818)) ;
    inv02 ix35167 (.Y (nx35168), .A (nx36820)) ;
    inv02 ix35169 (.Y (nx35170), .A (nx36820)) ;
    inv02 ix35171 (.Y (nx35172), .A (nx36820)) ;
    inv02 ix35173 (.Y (nx35174), .A (nx36820)) ;
    inv02 ix35175 (.Y (nx35176), .A (nx36820)) ;
    inv02 ix35177 (.Y (nx35178), .A (nx36820)) ;
    inv02 ix35179 (.Y (nx35180), .A (nx36820)) ;
    inv02 ix35181 (.Y (nx35182), .A (nx36822)) ;
    inv02 ix35183 (.Y (nx35184), .A (nx36822)) ;
    inv02 ix35185 (.Y (nx35186), .A (nx36822)) ;
    inv02 ix35187 (.Y (nx35188), .A (nx36822)) ;
    inv02 ix35189 (.Y (nx35190), .A (nx36822)) ;
    inv02 ix35191 (.Y (nx35192), .A (nx36822)) ;
    inv02 ix35193 (.Y (nx35194), .A (nx36822)) ;
    inv02 ix35195 (.Y (nx35196), .A (nx36824)) ;
    inv02 ix35197 (.Y (nx35198), .A (nx36824)) ;
    inv02 ix35199 (.Y (nx35200), .A (nx36824)) ;
    inv02 ix35201 (.Y (nx35202), .A (nx36824)) ;
    inv02 ix35203 (.Y (nx35204), .A (nx36824)) ;
    inv02 ix35205 (.Y (nx35206), .A (nx36824)) ;
    inv02 ix35207 (.Y (nx35208), .A (nx36824)) ;
    inv02 ix35209 (.Y (nx35210), .A (nx36826)) ;
    inv02 ix35211 (.Y (nx35212), .A (nx36826)) ;
    inv02 ix35215 (.Y (nx35216), .A (nx36828)) ;
    inv02 ix35217 (.Y (nx35218), .A (nx36828)) ;
    inv02 ix35219 (.Y (nx35220), .A (nx36828)) ;
    inv02 ix35221 (.Y (nx35222), .A (nx36828)) ;
    inv02 ix35223 (.Y (nx35224), .A (nx36828)) ;
    inv02 ix35225 (.Y (nx35226), .A (nx36828)) ;
    inv02 ix35227 (.Y (nx35228), .A (nx36828)) ;
    inv02 ix35229 (.Y (nx35230), .A (nx36830)) ;
    inv02 ix35231 (.Y (nx35232), .A (nx36830)) ;
    inv02 ix35233 (.Y (nx35234), .A (nx36830)) ;
    inv02 ix35235 (.Y (nx35236), .A (nx36830)) ;
    inv02 ix35237 (.Y (nx35238), .A (nx36830)) ;
    inv02 ix35239 (.Y (nx35240), .A (nx36830)) ;
    inv02 ix35241 (.Y (nx35242), .A (nx36830)) ;
    inv02 ix35243 (.Y (nx35244), .A (nx36832)) ;
    inv02 ix35245 (.Y (nx35246), .A (nx36832)) ;
    inv02 ix35247 (.Y (nx35248), .A (nx36832)) ;
    inv02 ix35249 (.Y (nx35250), .A (nx36832)) ;
    inv02 ix35251 (.Y (nx35252), .A (nx36832)) ;
    inv02 ix35253 (.Y (nx35254), .A (nx36832)) ;
    inv02 ix35255 (.Y (nx35256), .A (nx36832)) ;
    inv02 ix35257 (.Y (nx35258), .A (nx36834)) ;
    inv02 ix35259 (.Y (nx35260), .A (nx36834)) ;
    inv02 ix35261 (.Y (nx35262), .A (nx36834)) ;
    inv02 ix35263 (.Y (nx35264), .A (nx36834)) ;
    inv02 ix35265 (.Y (nx35266), .A (nx36834)) ;
    inv02 ix35267 (.Y (nx35268), .A (nx36834)) ;
    inv02 ix35269 (.Y (nx35270), .A (nx36834)) ;
    inv02 ix35271 (.Y (nx35272), .A (nx36836)) ;
    inv02 ix35273 (.Y (nx35274), .A (nx36836)) ;
    inv02 ix35275 (.Y (nx35276), .A (nx36836)) ;
    inv02 ix35277 (.Y (nx35278), .A (nx36836)) ;
    inv02 ix35279 (.Y (nx35280), .A (nx36836)) ;
    inv02 ix35281 (.Y (nx35282), .A (nx36836)) ;
    inv02 ix35283 (.Y (nx35284), .A (nx36836)) ;
    inv02 ix35285 (.Y (nx35286), .A (nx36838)) ;
    inv02 ix35287 (.Y (nx35288), .A (nx36838)) ;
    inv02 ix35291 (.Y (nx35292), .A (nx36840)) ;
    inv02 ix35293 (.Y (nx35294), .A (nx36840)) ;
    inv02 ix35295 (.Y (nx35296), .A (nx36840)) ;
    inv02 ix35297 (.Y (nx35298), .A (nx36840)) ;
    inv02 ix35299 (.Y (nx35300), .A (nx36840)) ;
    inv02 ix35301 (.Y (nx35302), .A (nx36840)) ;
    inv02 ix35303 (.Y (nx35304), .A (nx36840)) ;
    inv02 ix35305 (.Y (nx35306), .A (nx36842)) ;
    inv02 ix35307 (.Y (nx35308), .A (nx36842)) ;
    inv02 ix35309 (.Y (nx35310), .A (nx36842)) ;
    inv02 ix35311 (.Y (nx35312), .A (nx36842)) ;
    inv02 ix35313 (.Y (nx35314), .A (nx36842)) ;
    inv02 ix35315 (.Y (nx35316), .A (nx36842)) ;
    inv02 ix35317 (.Y (nx35318), .A (nx36842)) ;
    inv02 ix35319 (.Y (nx35320), .A (nx36844)) ;
    inv02 ix35321 (.Y (nx35322), .A (nx36844)) ;
    inv02 ix35323 (.Y (nx35324), .A (nx36844)) ;
    inv02 ix35325 (.Y (nx35326), .A (nx36844)) ;
    inv02 ix35327 (.Y (nx35328), .A (nx36844)) ;
    inv02 ix35329 (.Y (nx35330), .A (nx36844)) ;
    inv02 ix35331 (.Y (nx35332), .A (nx36844)) ;
    inv02 ix35333 (.Y (nx35334), .A (nx36846)) ;
    inv02 ix35335 (.Y (nx35336), .A (nx36846)) ;
    inv02 ix35337 (.Y (nx35338), .A (nx36846)) ;
    inv02 ix35339 (.Y (nx35340), .A (nx36846)) ;
    inv02 ix35341 (.Y (nx35342), .A (nx36846)) ;
    inv02 ix35343 (.Y (nx35344), .A (nx36846)) ;
    inv02 ix35345 (.Y (nx35346), .A (nx36846)) ;
    inv02 ix35347 (.Y (nx35348), .A (nx36848)) ;
    inv02 ix35349 (.Y (nx35350), .A (nx36848)) ;
    inv02 ix35351 (.Y (nx35352), .A (nx36848)) ;
    inv02 ix35353 (.Y (nx35354), .A (nx36848)) ;
    inv02 ix35355 (.Y (nx35356), .A (nx36848)) ;
    inv02 ix35357 (.Y (nx35358), .A (nx36848)) ;
    inv02 ix35359 (.Y (nx35360), .A (nx36848)) ;
    inv02 ix35361 (.Y (nx35362), .A (nx36850)) ;
    inv02 ix35363 (.Y (nx35364), .A (nx36850)) ;
    inv02 ix35367 (.Y (nx35368), .A (nx36852)) ;
    inv02 ix35369 (.Y (nx35370), .A (nx36852)) ;
    inv02 ix35371 (.Y (nx35372), .A (nx36852)) ;
    inv02 ix35373 (.Y (nx35374), .A (nx36852)) ;
    inv02 ix35375 (.Y (nx35376), .A (nx36852)) ;
    inv02 ix35377 (.Y (nx35378), .A (nx36852)) ;
    inv02 ix35379 (.Y (nx35380), .A (nx36852)) ;
    inv02 ix35381 (.Y (nx35382), .A (nx36854)) ;
    inv02 ix35383 (.Y (nx35384), .A (nx36854)) ;
    inv02 ix35385 (.Y (nx35386), .A (nx36854)) ;
    inv02 ix35387 (.Y (nx35388), .A (nx36854)) ;
    inv02 ix35389 (.Y (nx35390), .A (nx36854)) ;
    inv02 ix35391 (.Y (nx35392), .A (nx36854)) ;
    inv02 ix35393 (.Y (nx35394), .A (nx36854)) ;
    inv02 ix35395 (.Y (nx35396), .A (nx36856)) ;
    inv02 ix35397 (.Y (nx35398), .A (nx36856)) ;
    inv02 ix35399 (.Y (nx35400), .A (nx36856)) ;
    inv02 ix35401 (.Y (nx35402), .A (nx36856)) ;
    inv02 ix35403 (.Y (nx35404), .A (nx36856)) ;
    inv02 ix35405 (.Y (nx35406), .A (nx36856)) ;
    inv02 ix35407 (.Y (nx35408), .A (nx36856)) ;
    inv02 ix35409 (.Y (nx35410), .A (nx36858)) ;
    inv02 ix35411 (.Y (nx35412), .A (nx36858)) ;
    inv02 ix35413 (.Y (nx35414), .A (nx36858)) ;
    inv02 ix35415 (.Y (nx35416), .A (nx36858)) ;
    inv02 ix35417 (.Y (nx35418), .A (nx36858)) ;
    inv02 ix35419 (.Y (nx35420), .A (nx36858)) ;
    inv02 ix35421 (.Y (nx35422), .A (nx36858)) ;
    inv02 ix35423 (.Y (nx35424), .A (nx36860)) ;
    inv02 ix35425 (.Y (nx35426), .A (nx36860)) ;
    inv02 ix35427 (.Y (nx35428), .A (nx36860)) ;
    inv02 ix35429 (.Y (nx35430), .A (nx36860)) ;
    inv02 ix35431 (.Y (nx35432), .A (nx36860)) ;
    inv02 ix35433 (.Y (nx35434), .A (nx36860)) ;
    inv02 ix35435 (.Y (nx35436), .A (nx36860)) ;
    inv02 ix35437 (.Y (nx35438), .A (nx36862)) ;
    inv02 ix35439 (.Y (nx35440), .A (nx36862)) ;
    inv02 ix35443 (.Y (nx35444), .A (nx36864)) ;
    inv02 ix35445 (.Y (nx35446), .A (nx36864)) ;
    inv02 ix35447 (.Y (nx35448), .A (nx36864)) ;
    inv02 ix35449 (.Y (nx35450), .A (nx36864)) ;
    inv02 ix35451 (.Y (nx35452), .A (nx36864)) ;
    inv02 ix35453 (.Y (nx35454), .A (nx36864)) ;
    inv02 ix35455 (.Y (nx35456), .A (nx36864)) ;
    inv02 ix35457 (.Y (nx35458), .A (nx36866)) ;
    inv02 ix35459 (.Y (nx35460), .A (nx36866)) ;
    inv02 ix35461 (.Y (nx35462), .A (nx36866)) ;
    inv02 ix35463 (.Y (nx35464), .A (nx36866)) ;
    inv02 ix35465 (.Y (nx35466), .A (nx36866)) ;
    inv02 ix35467 (.Y (nx35468), .A (nx36866)) ;
    inv02 ix35469 (.Y (nx35470), .A (nx36866)) ;
    inv02 ix35471 (.Y (nx35472), .A (nx36868)) ;
    inv02 ix35473 (.Y (nx35474), .A (nx36868)) ;
    inv02 ix35475 (.Y (nx35476), .A (nx36868)) ;
    inv02 ix35477 (.Y (nx35478), .A (nx36868)) ;
    inv02 ix35479 (.Y (nx35480), .A (nx36868)) ;
    inv02 ix35481 (.Y (nx35482), .A (nx36868)) ;
    inv02 ix35483 (.Y (nx35484), .A (nx36868)) ;
    inv02 ix35485 (.Y (nx35486), .A (nx36870)) ;
    inv02 ix35487 (.Y (nx35488), .A (nx36870)) ;
    inv02 ix35489 (.Y (nx35490), .A (nx36870)) ;
    inv02 ix35491 (.Y (nx35492), .A (nx36870)) ;
    inv02 ix35493 (.Y (nx35494), .A (nx36870)) ;
    inv02 ix35495 (.Y (nx35496), .A (nx36870)) ;
    inv02 ix35497 (.Y (nx35498), .A (nx36870)) ;
    inv02 ix35499 (.Y (nx35500), .A (nx36872)) ;
    inv02 ix35501 (.Y (nx35502), .A (nx36872)) ;
    inv02 ix35503 (.Y (nx35504), .A (nx36872)) ;
    inv02 ix35505 (.Y (nx35506), .A (nx36872)) ;
    inv02 ix35507 (.Y (nx35508), .A (nx36872)) ;
    inv02 ix35509 (.Y (nx35510), .A (nx36872)) ;
    inv02 ix35511 (.Y (nx35512), .A (nx36872)) ;
    inv02 ix35513 (.Y (nx35514), .A (nx36874)) ;
    inv02 ix35515 (.Y (nx35516), .A (nx36874)) ;
    inv02 ix35519 (.Y (nx35520), .A (nx36876)) ;
    inv02 ix35521 (.Y (nx35522), .A (nx36876)) ;
    inv02 ix35523 (.Y (nx35524), .A (nx36876)) ;
    inv02 ix35525 (.Y (nx35526), .A (nx36876)) ;
    inv02 ix35527 (.Y (nx35528), .A (nx36876)) ;
    inv02 ix35529 (.Y (nx35530), .A (nx36876)) ;
    inv02 ix35531 (.Y (nx35532), .A (nx36876)) ;
    inv02 ix35533 (.Y (nx35534), .A (nx36878)) ;
    inv02 ix35535 (.Y (nx35536), .A (nx36878)) ;
    inv02 ix35537 (.Y (nx35538), .A (nx36878)) ;
    inv02 ix35539 (.Y (nx35540), .A (nx36878)) ;
    inv02 ix35541 (.Y (nx35542), .A (nx36878)) ;
    inv02 ix35543 (.Y (nx35544), .A (nx36878)) ;
    inv02 ix35545 (.Y (nx35546), .A (nx36878)) ;
    inv02 ix35547 (.Y (nx35548), .A (nx36880)) ;
    inv02 ix35549 (.Y (nx35550), .A (nx36880)) ;
    inv02 ix35551 (.Y (nx35552), .A (nx36880)) ;
    inv02 ix35553 (.Y (nx35554), .A (nx36880)) ;
    inv02 ix35555 (.Y (nx35556), .A (nx36880)) ;
    inv02 ix35557 (.Y (nx35558), .A (nx36880)) ;
    inv02 ix35559 (.Y (nx35560), .A (nx36880)) ;
    inv02 ix35561 (.Y (nx35562), .A (nx36882)) ;
    inv02 ix35563 (.Y (nx35564), .A (nx36882)) ;
    inv02 ix35565 (.Y (nx35566), .A (nx36882)) ;
    inv02 ix35567 (.Y (nx35568), .A (nx36882)) ;
    inv02 ix35569 (.Y (nx35570), .A (nx36882)) ;
    inv02 ix35571 (.Y (nx35572), .A (nx36882)) ;
    inv02 ix35573 (.Y (nx35574), .A (nx36882)) ;
    inv02 ix35575 (.Y (nx35576), .A (nx36884)) ;
    inv02 ix35577 (.Y (nx35578), .A (nx36884)) ;
    inv02 ix35579 (.Y (nx35580), .A (nx36884)) ;
    inv02 ix35581 (.Y (nx35582), .A (nx36884)) ;
    inv02 ix35583 (.Y (nx35584), .A (nx36884)) ;
    inv02 ix35585 (.Y (nx35586), .A (nx36884)) ;
    inv02 ix35587 (.Y (nx35588), .A (nx36884)) ;
    inv02 ix35589 (.Y (nx35590), .A (nx36886)) ;
    inv02 ix35591 (.Y (nx35592), .A (nx36886)) ;
    inv02 ix35595 (.Y (nx35596), .A (nx36888)) ;
    inv02 ix35597 (.Y (nx35598), .A (nx36888)) ;
    inv02 ix35599 (.Y (nx35600), .A (nx36888)) ;
    inv02 ix35601 (.Y (nx35602), .A (nx36888)) ;
    inv02 ix35603 (.Y (nx35604), .A (nx36888)) ;
    inv02 ix35605 (.Y (nx35606), .A (nx36888)) ;
    inv02 ix35607 (.Y (nx35608), .A (nx36888)) ;
    inv02 ix35609 (.Y (nx35610), .A (nx36890)) ;
    inv02 ix35611 (.Y (nx35612), .A (nx36890)) ;
    inv02 ix35613 (.Y (nx35614), .A (nx36890)) ;
    inv02 ix35615 (.Y (nx35616), .A (nx36890)) ;
    inv02 ix35617 (.Y (nx35618), .A (nx36890)) ;
    inv02 ix35619 (.Y (nx35620), .A (nx36890)) ;
    inv02 ix35621 (.Y (nx35622), .A (nx36890)) ;
    inv02 ix35623 (.Y (nx35624), .A (nx36892)) ;
    inv02 ix35625 (.Y (nx35626), .A (nx36892)) ;
    inv02 ix35627 (.Y (nx35628), .A (nx36892)) ;
    inv02 ix35629 (.Y (nx35630), .A (nx36892)) ;
    inv02 ix35631 (.Y (nx35632), .A (nx36892)) ;
    inv02 ix35633 (.Y (nx35634), .A (nx36892)) ;
    inv02 ix35635 (.Y (nx35636), .A (nx36892)) ;
    inv02 ix35637 (.Y (nx35638), .A (nx36894)) ;
    inv02 ix35639 (.Y (nx35640), .A (nx36894)) ;
    inv02 ix35641 (.Y (nx35642), .A (nx36894)) ;
    inv02 ix35643 (.Y (nx35644), .A (nx36894)) ;
    inv02 ix35645 (.Y (nx35646), .A (nx36894)) ;
    inv02 ix35647 (.Y (nx35648), .A (nx36894)) ;
    inv02 ix35649 (.Y (nx35650), .A (nx36894)) ;
    inv02 ix35651 (.Y (nx35652), .A (nx36896)) ;
    inv02 ix35653 (.Y (nx35654), .A (nx36896)) ;
    inv02 ix35655 (.Y (nx35656), .A (nx36896)) ;
    inv02 ix35657 (.Y (nx35658), .A (nx36896)) ;
    inv02 ix35659 (.Y (nx35660), .A (nx36896)) ;
    inv02 ix35661 (.Y (nx35662), .A (nx36896)) ;
    inv02 ix35663 (.Y (nx35664), .A (nx36896)) ;
    inv02 ix35665 (.Y (nx35666), .A (nx36898)) ;
    inv02 ix35667 (.Y (nx35668), .A (nx36898)) ;
    inv02 ix35669 (.Y (nx35670), .A (zero)) ;
    inv02 ix35671 (.Y (nx35672), .A (zero)) ;
    inv02 ix35673 (.Y (nx35674), .A (zero)) ;
    inv02 ix35675 (.Y (nx35676), .A (zero)) ;
    inv02 ix35677 (.Y (nx35678), .A (zero)) ;
    inv02 ix35679 (.Y (nx35680), .A (zero)) ;
    inv02 ix35681 (.Y (nx35682), .A (zero)) ;
    inv02 ix35683 (.Y (nx35684), .A (zero)) ;
    inv02 ix35685 (.Y (nx35686), .A (camera_module_algo_module_regs_rst)) ;
    inv02 ix35687 (.Y (nx35688), .A (nx37416)) ;
    inv02 ix35689 (.Y (nx35690), .A (nx37416)) ;
    inv02 ix35691 (.Y (nx35692), .A (rst)) ;
    inv02 ix35693 (.Y (nx35694), .A (rst)) ;
    inv02 ix35695 (.Y (nx35696), .A (nx879)) ;
    inv02 ix35697 (.Y (nx35698), .A (nx879)) ;
    inv02 ix35699 (.Y (nx35700), .A (nx25432)) ;
    inv02 ix35701 (.Y (nx35702), .A (nx37090)) ;
    inv02 ix35703 (.Y (nx35704), .A (nx37090)) ;
    inv02 ix35707 (.Y (nx35708), .A (nx37086)) ;
    buf02 ix35711 (.Y (nx35712), .A (nx22766)) ;
    buf02 ix35713 (.Y (nx35714), .A (nx22766)) ;
    inv02 ix35717 (.Y (nx35718), .A (camera_module_cache_address_from_DMA_0)) ;
    inv02 ix35719 (.Y (nx35720), .A (nx37412)) ;
    inv02 ix35781 (.Y (nx35782), .A (nx436)) ;
    inv02 ix35783 (.Y (nx35784), .A (nx436)) ;
    inv02 ix35785 (.Y (nx35786), .A (nx37370)) ;
    inv02 ix35795 (.Y (nx35796), .A (nx37074)) ;
    inv02 ix35803 (.Y (nx35804), .A (nx686)) ;
    inv02 ix35805 (.Y (nx35806), .A (nx686)) ;
    inv02 ix35807 (.Y (nx35808), .A (nx1490)) ;
    inv02 ix35809 (.Y (nx35810), .A (nx37404)) ;
    inv02 ix35811 (.Y (nx35812), .A (nx37404)) ;
    inv02 ix35813 (.Y (nx35814), .A (nx37404)) ;
    inv02 ix35815 (.Y (nx35816), .A (nx37404)) ;
    inv02 ix35817 (.Y (nx35818), .A (nx37404)) ;
    inv02 ix35819 (.Y (nx35820), .A (nx37404)) ;
    inv02 ix35821 (.Y (nx35822), .A (nx37404)) ;
    inv02 ix35823 (.Y (nx35824), .A (nx37010)) ;
    inv02 ix35825 (.Y (nx35826), .A (nx37010)) ;
    inv02 ix35827 (.Y (nx35828), .A (nx37010)) ;
    inv02 ix35829 (.Y (nx35830), .A (nx37010)) ;
    inv02 ix35831 (.Y (nx35832), .A (nx37010)) ;
    inv02 ix35833 (.Y (nx35834), .A (nx37010)) ;
    inv02 ix35835 (.Y (nx35836), .A (nx37010)) ;
    inv02 ix35837 (.Y (nx35838), .A (nx37012)) ;
    inv02 ix35839 (.Y (nx35840), .A (nx37012)) ;
    inv02 ix35841 (.Y (nx35842), .A (nx37012)) ;
    inv02 ix35843 (.Y (nx35844), .A (nx37012)) ;
    inv02 ix35845 (.Y (nx35846), .A (nx37012)) ;
    inv02 ix35847 (.Y (nx35848), .A (nx1472)) ;
    inv02 ix35849 (.Y (nx35850), .A (nx37402)) ;
    inv02 ix35851 (.Y (nx35852), .A (nx37402)) ;
    inv02 ix35853 (.Y (nx35854), .A (nx37402)) ;
    inv02 ix35855 (.Y (nx35856), .A (nx37402)) ;
    inv02 ix35857 (.Y (nx35858), .A (nx37402)) ;
    inv02 ix35859 (.Y (nx35860), .A (nx37402)) ;
    inv02 ix35861 (.Y (nx35862), .A (nx37402)) ;
    inv02 ix35863 (.Y (nx35864), .A (nx37004)) ;
    inv02 ix35865 (.Y (nx35866), .A (nx37004)) ;
    inv02 ix35867 (.Y (nx35868), .A (nx37004)) ;
    inv02 ix35869 (.Y (nx35870), .A (nx37004)) ;
    inv02 ix35871 (.Y (nx35872), .A (nx37004)) ;
    inv02 ix35873 (.Y (nx35874), .A (nx37004)) ;
    inv02 ix35875 (.Y (nx35876), .A (nx37004)) ;
    inv02 ix35877 (.Y (nx35878), .A (nx37006)) ;
    inv02 ix35879 (.Y (nx35880), .A (nx37006)) ;
    inv02 ix35881 (.Y (nx35882), .A (nx37006)) ;
    inv02 ix35883 (.Y (nx35884), .A (nx37006)) ;
    inv02 ix35885 (.Y (nx35886), .A (nx37006)) ;
    inv02 ix35887 (.Y (nx35888), .A (nx1452)) ;
    inv02 ix35889 (.Y (nx35890), .A (nx37400)) ;
    inv02 ix35891 (.Y (nx35892), .A (nx37400)) ;
    inv02 ix35893 (.Y (nx35894), .A (nx37400)) ;
    inv02 ix35895 (.Y (nx35896), .A (nx37400)) ;
    inv02 ix35897 (.Y (nx35898), .A (nx37400)) ;
    inv02 ix35899 (.Y (nx35900), .A (nx37400)) ;
    inv02 ix35901 (.Y (nx35902), .A (nx37400)) ;
    inv02 ix35903 (.Y (nx35904), .A (nx36998)) ;
    inv02 ix35905 (.Y (nx35906), .A (nx36998)) ;
    inv02 ix35907 (.Y (nx35908), .A (nx36998)) ;
    inv02 ix35909 (.Y (nx35910), .A (nx36998)) ;
    inv02 ix35911 (.Y (nx35912), .A (nx36998)) ;
    inv02 ix35913 (.Y (nx35914), .A (nx36998)) ;
    inv02 ix35915 (.Y (nx35916), .A (nx36998)) ;
    inv02 ix35917 (.Y (nx35918), .A (nx37000)) ;
    inv02 ix35919 (.Y (nx35920), .A (nx37000)) ;
    inv02 ix35921 (.Y (nx35922), .A (nx37000)) ;
    inv02 ix35923 (.Y (nx35924), .A (nx37000)) ;
    inv02 ix35925 (.Y (nx35926), .A (nx37000)) ;
    inv02 ix35927 (.Y (nx35928), .A (nx1434)) ;
    inv02 ix35929 (.Y (nx35930), .A (nx37398)) ;
    inv02 ix35931 (.Y (nx35932), .A (nx37398)) ;
    inv02 ix35933 (.Y (nx35934), .A (nx37398)) ;
    inv02 ix35935 (.Y (nx35936), .A (nx37398)) ;
    inv02 ix35937 (.Y (nx35938), .A (nx37398)) ;
    inv02 ix35939 (.Y (nx35940), .A (nx37398)) ;
    inv02 ix35941 (.Y (nx35942), .A (nx37398)) ;
    inv02 ix35943 (.Y (nx35944), .A (nx36992)) ;
    inv02 ix35945 (.Y (nx35946), .A (nx36992)) ;
    inv02 ix35947 (.Y (nx35948), .A (nx36992)) ;
    inv02 ix35949 (.Y (nx35950), .A (nx36992)) ;
    inv02 ix35951 (.Y (nx35952), .A (nx36992)) ;
    inv02 ix35953 (.Y (nx35954), .A (nx36992)) ;
    inv02 ix35955 (.Y (nx35956), .A (nx36992)) ;
    inv02 ix35957 (.Y (nx35958), .A (nx36994)) ;
    inv02 ix35959 (.Y (nx35960), .A (nx36994)) ;
    inv02 ix35961 (.Y (nx35962), .A (nx36994)) ;
    inv02 ix35963 (.Y (nx35964), .A (nx36994)) ;
    inv02 ix35965 (.Y (nx35966), .A (nx36994)) ;
    inv02 ix35967 (.Y (nx35968), .A (nx1410)) ;
    inv02 ix35969 (.Y (nx35970), .A (nx37396)) ;
    inv02 ix35971 (.Y (nx35972), .A (nx37396)) ;
    inv02 ix35973 (.Y (nx35974), .A (nx37396)) ;
    inv02 ix35975 (.Y (nx35976), .A (nx37396)) ;
    inv02 ix35977 (.Y (nx35978), .A (nx37396)) ;
    inv02 ix35979 (.Y (nx35980), .A (nx37396)) ;
    inv02 ix35981 (.Y (nx35982), .A (nx37396)) ;
    inv02 ix35983 (.Y (nx35984), .A (nx36986)) ;
    inv02 ix35985 (.Y (nx35986), .A (nx36986)) ;
    inv02 ix35987 (.Y (nx35988), .A (nx36986)) ;
    inv02 ix35989 (.Y (nx35990), .A (nx36986)) ;
    inv02 ix35991 (.Y (nx35992), .A (nx36986)) ;
    inv02 ix35993 (.Y (nx35994), .A (nx36986)) ;
    inv02 ix35995 (.Y (nx35996), .A (nx36986)) ;
    inv02 ix35997 (.Y (nx35998), .A (nx36988)) ;
    inv02 ix35999 (.Y (nx36000), .A (nx36988)) ;
    inv02 ix36001 (.Y (nx36002), .A (nx36988)) ;
    inv02 ix36003 (.Y (nx36004), .A (nx36988)) ;
    inv02 ix36005 (.Y (nx36006), .A (nx36988)) ;
    inv02 ix36007 (.Y (nx36008), .A (nx1392)) ;
    inv02 ix36009 (.Y (nx36010), .A (nx37394)) ;
    inv02 ix36011 (.Y (nx36012), .A (nx37394)) ;
    inv02 ix36013 (.Y (nx36014), .A (nx37394)) ;
    inv02 ix36015 (.Y (nx36016), .A (nx37394)) ;
    inv02 ix36017 (.Y (nx36018), .A (nx37394)) ;
    inv02 ix36019 (.Y (nx36020), .A (nx37394)) ;
    inv02 ix36021 (.Y (nx36022), .A (nx37394)) ;
    inv02 ix36023 (.Y (nx36024), .A (nx36980)) ;
    inv02 ix36025 (.Y (nx36026), .A (nx36980)) ;
    inv02 ix36027 (.Y (nx36028), .A (nx36980)) ;
    inv02 ix36029 (.Y (nx36030), .A (nx36980)) ;
    inv02 ix36031 (.Y (nx36032), .A (nx36980)) ;
    inv02 ix36033 (.Y (nx36034), .A (nx36980)) ;
    inv02 ix36035 (.Y (nx36036), .A (nx36980)) ;
    inv02 ix36037 (.Y (nx36038), .A (nx36982)) ;
    inv02 ix36039 (.Y (nx36040), .A (nx36982)) ;
    inv02 ix36041 (.Y (nx36042), .A (nx36982)) ;
    inv02 ix36043 (.Y (nx36044), .A (nx36982)) ;
    inv02 ix36045 (.Y (nx36046), .A (nx36982)) ;
    inv02 ix36047 (.Y (nx36048), .A (nx1354)) ;
    inv02 ix36049 (.Y (nx36050), .A (nx37390)) ;
    inv02 ix36051 (.Y (nx36052), .A (nx37390)) ;
    inv02 ix36053 (.Y (nx36054), .A (nx37390)) ;
    inv02 ix36055 (.Y (nx36056), .A (nx37390)) ;
    inv02 ix36057 (.Y (nx36058), .A (nx37390)) ;
    inv02 ix36059 (.Y (nx36060), .A (nx37390)) ;
    inv02 ix36061 (.Y (nx36062), .A (nx37390)) ;
    inv02 ix36063 (.Y (nx36064), .A (nx36968)) ;
    inv02 ix36065 (.Y (nx36066), .A (nx36968)) ;
    inv02 ix36067 (.Y (nx36068), .A (nx36968)) ;
    inv02 ix36069 (.Y (nx36070), .A (nx36968)) ;
    inv02 ix36071 (.Y (nx36072), .A (nx36968)) ;
    inv02 ix36073 (.Y (nx36074), .A (nx36968)) ;
    inv02 ix36075 (.Y (nx36076), .A (nx36968)) ;
    inv02 ix36077 (.Y (nx36078), .A (nx36970)) ;
    inv02 ix36079 (.Y (nx36080), .A (nx36970)) ;
    inv02 ix36081 (.Y (nx36082), .A (nx36970)) ;
    inv02 ix36083 (.Y (nx36084), .A (nx36970)) ;
    inv02 ix36085 (.Y (nx36086), .A (nx36970)) ;
    inv02 ix36087 (.Y (nx36088), .A (nx1372)) ;
    inv02 ix36089 (.Y (nx36090), .A (nx37392)) ;
    inv02 ix36091 (.Y (nx36092), .A (nx37392)) ;
    inv02 ix36093 (.Y (nx36094), .A (nx37392)) ;
    inv02 ix36095 (.Y (nx36096), .A (nx37392)) ;
    inv02 ix36097 (.Y (nx36098), .A (nx37392)) ;
    inv02 ix36099 (.Y (nx36100), .A (nx37392)) ;
    inv02 ix36101 (.Y (nx36102), .A (nx37392)) ;
    inv02 ix36103 (.Y (nx36104), .A (nx36974)) ;
    inv02 ix36105 (.Y (nx36106), .A (nx36974)) ;
    inv02 ix36107 (.Y (nx36108), .A (nx36974)) ;
    inv02 ix36109 (.Y (nx36110), .A (nx36974)) ;
    inv02 ix36111 (.Y (nx36112), .A (nx36974)) ;
    inv02 ix36113 (.Y (nx36114), .A (nx36974)) ;
    inv02 ix36115 (.Y (nx36116), .A (nx36974)) ;
    inv02 ix36117 (.Y (nx36118), .A (nx36976)) ;
    inv02 ix36119 (.Y (nx36120), .A (nx36976)) ;
    inv02 ix36121 (.Y (nx36122), .A (nx36976)) ;
    inv02 ix36123 (.Y (nx36124), .A (nx36976)) ;
    inv02 ix36125 (.Y (nx36126), .A (nx36976)) ;
    inv02 ix36127 (.Y (nx36128), .A (nx1326)) ;
    inv02 ix36129 (.Y (nx36130), .A (nx37388)) ;
    inv02 ix36131 (.Y (nx36132), .A (nx37388)) ;
    inv02 ix36133 (.Y (nx36134), .A (nx37388)) ;
    inv02 ix36135 (.Y (nx36136), .A (nx37388)) ;
    inv02 ix36137 (.Y (nx36138), .A (nx37388)) ;
    inv02 ix36139 (.Y (nx36140), .A (nx37388)) ;
    inv02 ix36141 (.Y (nx36142), .A (nx37388)) ;
    inv02 ix36143 (.Y (nx36144), .A (nx36962)) ;
    inv02 ix36145 (.Y (nx36146), .A (nx36962)) ;
    inv02 ix36147 (.Y (nx36148), .A (nx36962)) ;
    inv02 ix36149 (.Y (nx36150), .A (nx36962)) ;
    inv02 ix36151 (.Y (nx36152), .A (nx36962)) ;
    inv02 ix36153 (.Y (nx36154), .A (nx36962)) ;
    inv02 ix36155 (.Y (nx36156), .A (nx36962)) ;
    inv02 ix36157 (.Y (nx36158), .A (nx36964)) ;
    inv02 ix36159 (.Y (nx36160), .A (nx36964)) ;
    inv02 ix36161 (.Y (nx36162), .A (nx36964)) ;
    inv02 ix36163 (.Y (nx36164), .A (nx36964)) ;
    inv02 ix36165 (.Y (nx36166), .A (nx36964)) ;
    inv02 ix36167 (.Y (nx36168), .A (nx1308)) ;
    inv02 ix36169 (.Y (nx36170), .A (nx37386)) ;
    inv02 ix36171 (.Y (nx36172), .A (nx37386)) ;
    inv02 ix36173 (.Y (nx36174), .A (nx37386)) ;
    inv02 ix36175 (.Y (nx36176), .A (nx37386)) ;
    inv02 ix36177 (.Y (nx36178), .A (nx37386)) ;
    inv02 ix36179 (.Y (nx36180), .A (nx37386)) ;
    inv02 ix36181 (.Y (nx36182), .A (nx37386)) ;
    inv02 ix36183 (.Y (nx36184), .A (nx36956)) ;
    inv02 ix36185 (.Y (nx36186), .A (nx36956)) ;
    inv02 ix36187 (.Y (nx36188), .A (nx36956)) ;
    inv02 ix36189 (.Y (nx36190), .A (nx36956)) ;
    inv02 ix36191 (.Y (nx36192), .A (nx36956)) ;
    inv02 ix36193 (.Y (nx36194), .A (nx36956)) ;
    inv02 ix36195 (.Y (nx36196), .A (nx36956)) ;
    inv02 ix36197 (.Y (nx36198), .A (nx36958)) ;
    inv02 ix36199 (.Y (nx36200), .A (nx36958)) ;
    inv02 ix36201 (.Y (nx36202), .A (nx36958)) ;
    inv02 ix36203 (.Y (nx36204), .A (nx36958)) ;
    inv02 ix36205 (.Y (nx36206), .A (nx36958)) ;
    inv02 ix36207 (.Y (nx36208), .A (nx1270)) ;
    inv02 ix36209 (.Y (nx36210), .A (nx37382)) ;
    inv02 ix36211 (.Y (nx36212), .A (nx37382)) ;
    inv02 ix36213 (.Y (nx36214), .A (nx37382)) ;
    inv02 ix36215 (.Y (nx36216), .A (nx37382)) ;
    inv02 ix36217 (.Y (nx36218), .A (nx37382)) ;
    inv02 ix36219 (.Y (nx36220), .A (nx37382)) ;
    inv02 ix36221 (.Y (nx36222), .A (nx37382)) ;
    inv02 ix36223 (.Y (nx36224), .A (nx36944)) ;
    inv02 ix36225 (.Y (nx36226), .A (nx36944)) ;
    inv02 ix36227 (.Y (nx36228), .A (nx36944)) ;
    inv02 ix36229 (.Y (nx36230), .A (nx36944)) ;
    inv02 ix36231 (.Y (nx36232), .A (nx36944)) ;
    inv02 ix36233 (.Y (nx36234), .A (nx36944)) ;
    inv02 ix36235 (.Y (nx36236), .A (nx36944)) ;
    inv02 ix36237 (.Y (nx36238), .A (nx36946)) ;
    inv02 ix36239 (.Y (nx36240), .A (nx36946)) ;
    inv02 ix36241 (.Y (nx36242), .A (nx36946)) ;
    inv02 ix36243 (.Y (nx36244), .A (nx36946)) ;
    inv02 ix36245 (.Y (nx36246), .A (nx36946)) ;
    inv02 ix36247 (.Y (nx36248), .A (nx1288)) ;
    inv02 ix36249 (.Y (nx36250), .A (nx37384)) ;
    inv02 ix36251 (.Y (nx36252), .A (nx37384)) ;
    inv02 ix36253 (.Y (nx36254), .A (nx37384)) ;
    inv02 ix36255 (.Y (nx36256), .A (nx37384)) ;
    inv02 ix36257 (.Y (nx36258), .A (nx37384)) ;
    inv02 ix36259 (.Y (nx36260), .A (nx37384)) ;
    inv02 ix36261 (.Y (nx36262), .A (nx37384)) ;
    inv02 ix36263 (.Y (nx36264), .A (nx36950)) ;
    inv02 ix36265 (.Y (nx36266), .A (nx36950)) ;
    inv02 ix36267 (.Y (nx36268), .A (nx36950)) ;
    inv02 ix36269 (.Y (nx36270), .A (nx36950)) ;
    inv02 ix36271 (.Y (nx36272), .A (nx36950)) ;
    inv02 ix36273 (.Y (nx36274), .A (nx36950)) ;
    inv02 ix36275 (.Y (nx36276), .A (nx36950)) ;
    inv02 ix36277 (.Y (nx36278), .A (nx36952)) ;
    inv02 ix36279 (.Y (nx36280), .A (nx36952)) ;
    inv02 ix36281 (.Y (nx36282), .A (nx36952)) ;
    inv02 ix36283 (.Y (nx36284), .A (nx36952)) ;
    inv02 ix36285 (.Y (nx36286), .A (nx36952)) ;
    inv02 ix36287 (.Y (nx36288), .A (nx37380)) ;
    inv02 ix36289 (.Y (nx36290), .A (nx37380)) ;
    inv02 ix36291 (.Y (nx36292), .A (nx37380)) ;
    inv02 ix36293 (.Y (nx36294), .A (nx37380)) ;
    inv02 ix36295 (.Y (nx36296), .A (nx37380)) ;
    inv02 ix36297 (.Y (nx36298), .A (nx37380)) ;
    inv02 ix36299 (.Y (nx36300), .A (nx37380)) ;
    inv02 ix36301 (.Y (nx36302), .A (nx36938)) ;
    inv02 ix36303 (.Y (nx36304), .A (nx36938)) ;
    inv02 ix36305 (.Y (nx36306), .A (nx36938)) ;
    inv02 ix36307 (.Y (nx36308), .A (nx36938)) ;
    inv02 ix36309 (.Y (nx36310), .A (nx36938)) ;
    inv02 ix36311 (.Y (nx36312), .A (nx36938)) ;
    inv02 ix36313 (.Y (nx36314), .A (nx36938)) ;
    inv02 ix36315 (.Y (nx36316), .A (nx36940)) ;
    inv02 ix36317 (.Y (nx36318), .A (nx36940)) ;
    inv02 ix36319 (.Y (nx36320), .A (nx36940)) ;
    inv02 ix36321 (.Y (nx36322), .A (nx36940)) ;
    inv02 ix36323 (.Y (nx36324), .A (nx36940)) ;
    inv02 ix36325 (.Y (nx36326), .A (nx36940)) ;
    inv02 ix36327 (.Y (nx36328), .A (nx37378)) ;
    inv02 ix36329 (.Y (nx36330), .A (nx37378)) ;
    inv02 ix36331 (.Y (nx36332), .A (nx37378)) ;
    inv02 ix36333 (.Y (nx36334), .A (nx37378)) ;
    inv02 ix36335 (.Y (nx36336), .A (nx37378)) ;
    inv02 ix36337 (.Y (nx36338), .A (nx37378)) ;
    inv02 ix36339 (.Y (nx36340), .A (nx37378)) ;
    inv02 ix36341 (.Y (nx36342), .A (nx36932)) ;
    inv02 ix36343 (.Y (nx36344), .A (nx36932)) ;
    inv02 ix36345 (.Y (nx36346), .A (nx36932)) ;
    inv02 ix36347 (.Y (nx36348), .A (nx36932)) ;
    inv02 ix36349 (.Y (nx36350), .A (nx36932)) ;
    inv02 ix36351 (.Y (nx36352), .A (nx36932)) ;
    inv02 ix36353 (.Y (nx36354), .A (nx36932)) ;
    inv02 ix36355 (.Y (nx36356), .A (nx36934)) ;
    inv02 ix36357 (.Y (nx36358), .A (nx36934)) ;
    inv02 ix36359 (.Y (nx36360), .A (nx36934)) ;
    inv02 ix36361 (.Y (nx36362), .A (nx36934)) ;
    inv02 ix36363 (.Y (nx36364), .A (nx36934)) ;
    inv02 ix36365 (.Y (nx36366), .A (nx36934)) ;
    inv02 ix36367 (.Y (nx36368), .A (nx37376)) ;
    inv02 ix36369 (.Y (nx36370), .A (nx37376)) ;
    inv02 ix36371 (.Y (nx36372), .A (nx37376)) ;
    inv02 ix36373 (.Y (nx36374), .A (nx37376)) ;
    inv02 ix36375 (.Y (nx36376), .A (nx37376)) ;
    inv02 ix36377 (.Y (nx36378), .A (nx37376)) ;
    inv02 ix36379 (.Y (nx36380), .A (nx37376)) ;
    inv02 ix36381 (.Y (nx36382), .A (nx36926)) ;
    inv02 ix36383 (.Y (nx36384), .A (nx36926)) ;
    inv02 ix36385 (.Y (nx36386), .A (nx36926)) ;
    inv02 ix36387 (.Y (nx36388), .A (nx36926)) ;
    inv02 ix36389 (.Y (nx36390), .A (nx36926)) ;
    inv02 ix36391 (.Y (nx36392), .A (nx36926)) ;
    inv02 ix36393 (.Y (nx36394), .A (nx36926)) ;
    inv02 ix36395 (.Y (nx36396), .A (nx36928)) ;
    inv02 ix36397 (.Y (nx36398), .A (nx36928)) ;
    inv02 ix36399 (.Y (nx36400), .A (nx36928)) ;
    inv02 ix36401 (.Y (nx36402), .A (nx36928)) ;
    inv02 ix36403 (.Y (nx36404), .A (nx36928)) ;
    inv02 ix36405 (.Y (nx36406), .A (nx36928)) ;
    inv02 ix36407 (.Y (nx36408), .A (nx37374)) ;
    inv02 ix36409 (.Y (nx36410), .A (nx37374)) ;
    inv02 ix36411 (.Y (nx36412), .A (nx37374)) ;
    inv02 ix36413 (.Y (nx36414), .A (nx37374)) ;
    inv02 ix36415 (.Y (nx36416), .A (nx37374)) ;
    inv02 ix36417 (.Y (nx36418), .A (nx37374)) ;
    inv02 ix36419 (.Y (nx36420), .A (nx37374)) ;
    inv02 ix36421 (.Y (nx36422), .A (nx36918)) ;
    inv02 ix36423 (.Y (nx36424), .A (nx36918)) ;
    inv02 ix36425 (.Y (nx36426), .A (nx36918)) ;
    inv02 ix36427 (.Y (nx36428), .A (nx36918)) ;
    inv02 ix36429 (.Y (nx36430), .A (nx36918)) ;
    inv02 ix36431 (.Y (nx36432), .A (nx36918)) ;
    inv02 ix36433 (.Y (nx36434), .A (nx36918)) ;
    inv02 ix36435 (.Y (nx36436), .A (nx36920)) ;
    inv02 ix36437 (.Y (nx36438), .A (nx36920)) ;
    inv02 ix36439 (.Y (nx36440), .A (nx36920)) ;
    inv02 ix36441 (.Y (nx36442), .A (nx36920)) ;
    inv02 ix36443 (.Y (nx36444), .A (nx36920)) ;
    inv02 ix36445 (.Y (nx36446), .A (nx36920)) ;
    inv02 ix36447 (.Y (nx36448), .A (nx5650)) ;
    inv02 ix36449 (.Y (nx36450), .A (nx5650)) ;
    inv02 ix36451 (.Y (nx36452), .A (nx5358)) ;
    inv02 ix36453 (.Y (nx36454), .A (nx5358)) ;
    inv02 ix36455 (.Y (nx36456), .A (nx5064)) ;
    inv02 ix36457 (.Y (nx36458), .A (nx5064)) ;
    inv02 ix36459 (.Y (nx36460), .A (nx4772)) ;
    inv02 ix36461 (.Y (nx36462), .A (nx4772)) ;
    inv02 ix36463 (.Y (nx36464), .A (nx4474)) ;
    inv02 ix36465 (.Y (nx36466), .A (nx4474)) ;
    inv02 ix36467 (.Y (nx36468), .A (nx4182)) ;
    inv02 ix36469 (.Y (nx36470), .A (nx4182)) ;
    inv02 ix36471 (.Y (nx36472), .A (nx3888)) ;
    inv02 ix36473 (.Y (nx36474), .A (nx3888)) ;
    inv02 ix36475 (.Y (nx36476), .A (nx3596)) ;
    inv02 ix36477 (.Y (nx36478), .A (nx3596)) ;
    inv02 ix36479 (.Y (nx36480), .A (nx3294)) ;
    inv02 ix36481 (.Y (nx36482), .A (nx3294)) ;
    inv02 ix36483 (.Y (nx36484), .A (nx3002)) ;
    inv02 ix36485 (.Y (nx36486), .A (nx3002)) ;
    inv02 ix36487 (.Y (nx36488), .A (nx2708)) ;
    inv02 ix36489 (.Y (nx36490), .A (nx2708)) ;
    inv02 ix36491 (.Y (nx36492), .A (nx2416)) ;
    inv02 ix36493 (.Y (nx36494), .A (nx2416)) ;
    buf02 ix36495 (.Y (nx36496), .A (nx24463)) ;
    buf02 ix36497 (.Y (nx36498), .A (nx24463)) ;
    inv02 ix36505 (.Y (nx36506), .A (nx36500)) ;
    inv02 ix36507 (.Y (nx36508), .A (nx37280)) ;
    buf02 ix36509 (.Y (nx36510), .A (nx24473)) ;
    buf02 ix36511 (.Y (nx36512), .A (nx24473)) ;
    buf02 ix36513 (.Y (nx36514), .A (nx24481)) ;
    buf02 ix36515 (.Y (nx36516), .A (nx24481)) ;
    buf02 ix36517 (.Y (nx36518), .A (nx24487)) ;
    buf02 ix36519 (.Y (nx36520), .A (nx24487)) ;
    buf02 ix36521 (.Y (nx36522), .A (nx24495)) ;
    buf02 ix36523 (.Y (nx36524), .A (nx24495)) ;
    buf02 ix36525 (.Y (nx36526), .A (nx24500)) ;
    buf02 ix36527 (.Y (nx36528), .A (nx24500)) ;
    buf02 ix36529 (.Y (nx36530), .A (nx24508)) ;
    buf02 ix36531 (.Y (nx36532), .A (nx24508)) ;
    buf02 ix36533 (.Y (nx36534), .A (nx24513)) ;
    buf02 ix36535 (.Y (nx36536), .A (nx24513)) ;
    buf02 ix36537 (.Y (nx36538), .A (nx24521)) ;
    buf02 ix36539 (.Y (nx36540), .A (nx24521)) ;
    buf02 ix36541 (.Y (nx36542), .A (nx24526)) ;
    buf02 ix36543 (.Y (nx36544), .A (nx24526)) ;
    buf02 ix36545 (.Y (nx36546), .A (nx24535)) ;
    buf02 ix36547 (.Y (nx36548), .A (nx24535)) ;
    buf02 ix36549 (.Y (nx36550), .A (nx24541)) ;
    buf02 ix36551 (.Y (nx36552), .A (nx24541)) ;
    buf02 ix36553 (.Y (nx36554), .A (nx24548)) ;
    buf02 ix36555 (.Y (nx36556), .A (nx24548)) ;
    buf02 ix36557 (.Y (nx36558), .A (nx24554)) ;
    buf02 ix36559 (.Y (nx36560), .A (nx24554)) ;
    buf02 ix36561 (.Y (nx36562), .A (nx24563)) ;
    buf02 ix36563 (.Y (nx36564), .A (nx24563)) ;
    buf02 ix36565 (.Y (nx36566), .A (nx24569)) ;
    buf02 ix36567 (.Y (nx36568), .A (nx24569)) ;
    buf02 ix36569 (.Y (nx36570), .A (nx24581)) ;
    buf02 ix36571 (.Y (nx36572), .A (nx24581)) ;
    inv02 ix36579 (.Y (nx36580), .A (nx36574)) ;
    inv02 ix36581 (.Y (nx36582), .A (nx37286)) ;
    buf02 ix36583 (.Y (nx36584), .A (nx24589)) ;
    buf02 ix36585 (.Y (nx36586), .A (nx24589)) ;
    buf02 ix36587 (.Y (nx36588), .A (nx24597)) ;
    buf02 ix36589 (.Y (nx36590), .A (nx24597)) ;
    buf02 ix36591 (.Y (nx36592), .A (nx24602)) ;
    buf02 ix36593 (.Y (nx36594), .A (nx24602)) ;
    buf02 ix36595 (.Y (nx36596), .A (nx24610)) ;
    buf02 ix36597 (.Y (nx36598), .A (nx24610)) ;
    buf02 ix36599 (.Y (nx36600), .A (nx24615)) ;
    buf02 ix36601 (.Y (nx36602), .A (nx24615)) ;
    buf02 ix36603 (.Y (nx36604), .A (nx24624)) ;
    buf02 ix36605 (.Y (nx36606), .A (nx24624)) ;
    buf02 ix36607 (.Y (nx36608), .A (nx24629)) ;
    buf02 ix36609 (.Y (nx36610), .A (nx24629)) ;
    buf02 ix36611 (.Y (nx36612), .A (nx24637)) ;
    buf02 ix36613 (.Y (nx36614), .A (nx24637)) ;
    buf02 ix36615 (.Y (nx36616), .A (nx24642)) ;
    buf02 ix36617 (.Y (nx36618), .A (nx24642)) ;
    buf02 ix36619 (.Y (nx36620), .A (nx24650)) ;
    buf02 ix36621 (.Y (nx36622), .A (nx24650)) ;
    buf02 ix36623 (.Y (nx36624), .A (nx24655)) ;
    buf02 ix36625 (.Y (nx36626), .A (nx24655)) ;
    buf02 ix36627 (.Y (nx36628), .A (nx24663)) ;
    buf02 ix36629 (.Y (nx36630), .A (nx24663)) ;
    buf02 ix36631 (.Y (nx36632), .A (nx24669)) ;
    buf02 ix36633 (.Y (nx36634), .A (nx24669)) ;
    buf02 ix36635 (.Y (nx36636), .A (nx24677)) ;
    buf02 ix36637 (.Y (nx36638), .A (nx24677)) ;
    buf02 ix36639 (.Y (nx36640), .A (nx24682)) ;
    buf02 ix36641 (.Y (nx36642), .A (nx24682)) ;
    buf02 ix36643 (.Y (nx36644), .A (nx24693)) ;
    buf02 ix36645 (.Y (nx36646), .A (nx24693)) ;
    inv02 ix36653 (.Y (nx36654), .A (nx36648)) ;
    inv02 ix36655 (.Y (nx36656), .A (nx37292)) ;
    buf02 ix36657 (.Y (nx36658), .A (nx24703)) ;
    buf02 ix36659 (.Y (nx36660), .A (nx24703)) ;
    buf02 ix36661 (.Y (nx36662), .A (nx24712)) ;
    buf02 ix36663 (.Y (nx36664), .A (nx24712)) ;
    buf02 ix36665 (.Y (nx36666), .A (nx24717)) ;
    buf02 ix36667 (.Y (nx36668), .A (nx24717)) ;
    buf02 ix36669 (.Y (nx36670), .A (nx24725)) ;
    buf02 ix36671 (.Y (nx36672), .A (nx24725)) ;
    buf02 ix36673 (.Y (nx36674), .A (nx24730)) ;
    buf02 ix36675 (.Y (nx36676), .A (nx24730)) ;
    buf02 ix36677 (.Y (nx36678), .A (nx24738)) ;
    buf02 ix36679 (.Y (nx36680), .A (nx24738)) ;
    buf02 ix36681 (.Y (nx36682), .A (nx24743)) ;
    buf02 ix36683 (.Y (nx36684), .A (nx24743)) ;
    buf02 ix36685 (.Y (nx36686), .A (nx24751)) ;
    buf02 ix36687 (.Y (nx36688), .A (nx24751)) ;
    buf02 ix36689 (.Y (nx36690), .A (nx24757)) ;
    buf02 ix36691 (.Y (nx36692), .A (nx24757)) ;
    buf02 ix36693 (.Y (nx36694), .A (nx24765)) ;
    buf02 ix36695 (.Y (nx36696), .A (nx24765)) ;
    buf02 ix36697 (.Y (nx36698), .A (nx24770)) ;
    buf02 ix36699 (.Y (nx36700), .A (nx24770)) ;
    buf02 ix36701 (.Y (nx36702), .A (nx24778)) ;
    buf02 ix36703 (.Y (nx36704), .A (nx24778)) ;
    buf02 ix36705 (.Y (nx36706), .A (nx24785)) ;
    buf02 ix36707 (.Y (nx36708), .A (nx24785)) ;
    buf02 ix36709 (.Y (nx36710), .A (nx24792)) ;
    buf02 ix36711 (.Y (nx36712), .A (nx24792)) ;
    buf02 ix36713 (.Y (nx36714), .A (nx24798)) ;
    buf02 ix36715 (.Y (nx36716), .A (nx24798)) ;
    buf02 ix36717 (.Y (nx36718), .A (nx24809)) ;
    buf02 ix36719 (.Y (nx36720), .A (nx24809)) ;
    inv02 ix36727 (.Y (nx36728), .A (nx37298)) ;
    inv02 ix36729 (.Y (nx36730), .A (nx37298)) ;
    buf02 ix36731 (.Y (nx36732), .A (nx24816)) ;
    buf02 ix36733 (.Y (nx36734), .A (nx24816)) ;
    buf02 ix36735 (.Y (nx36736), .A (nx24825)) ;
    buf02 ix36737 (.Y (nx36738), .A (nx24825)) ;
    buf02 ix36739 (.Y (nx36740), .A (nx24830)) ;
    buf02 ix36741 (.Y (nx36742), .A (nx24830)) ;
    buf02 ix36743 (.Y (nx36744), .A (nx24838)) ;
    buf02 ix36745 (.Y (nx36746), .A (nx24838)) ;
    buf02 ix36747 (.Y (nx36748), .A (nx24845)) ;
    buf02 ix36749 (.Y (nx36750), .A (nx24845)) ;
    buf02 ix36751 (.Y (nx36752), .A (nx24853)) ;
    buf02 ix36753 (.Y (nx36754), .A (nx24853)) ;
    buf02 ix36755 (.Y (nx36756), .A (nx24859)) ;
    buf02 ix36757 (.Y (nx36758), .A (nx24859)) ;
    buf02 ix36759 (.Y (nx36760), .A (nx24869)) ;
    buf02 ix36761 (.Y (nx36762), .A (nx24869)) ;
    buf02 ix36763 (.Y (nx36764), .A (nx24874)) ;
    buf02 ix36765 (.Y (nx36766), .A (nx24874)) ;
    buf02 ix36767 (.Y (nx36768), .A (nx24882)) ;
    buf02 ix36769 (.Y (nx36770), .A (nx24882)) ;
    buf02 ix36771 (.Y (nx36772), .A (nx24887)) ;
    buf02 ix36773 (.Y (nx36774), .A (nx24887)) ;
    buf02 ix36775 (.Y (nx36776), .A (nx24894)) ;
    buf02 ix36777 (.Y (nx36778), .A (nx24894)) ;
    buf02 ix36779 (.Y (nx36780), .A (nx24900)) ;
    buf02 ix36781 (.Y (nx36782), .A (nx24900)) ;
    buf02 ix36783 (.Y (nx36784), .A (nx24909)) ;
    buf02 ix36785 (.Y (nx36786), .A (nx24909)) ;
    buf02 ix36787 (.Y (nx36788), .A (nx24914)) ;
    buf02 ix36789 (.Y (nx36790), .A (nx24914)) ;
    buf02 ix36791 (.Y (nx36792), .A (nx24918)) ;
    buf02 ix36793 (.Y (nx36794), .A (nx24918)) ;
    inv02 ix36803 (.Y (nx36804), .A (nx1186)) ;
    inv02 ix36805 (.Y (nx36806), .A (nx36922)) ;
    inv02 ix36807 (.Y (nx36808), .A (nx36922)) ;
    inv02 ix36809 (.Y (nx36810), .A (nx36922)) ;
    inv02 ix36811 (.Y (nx36812), .A (nx36922)) ;
    inv02 ix36813 (.Y (nx36814), .A (nx36922)) ;
    inv02 ix36815 (.Y (nx36816), .A (nx6100)) ;
    inv02 ix36817 (.Y (nx36818), .A (nx37014)) ;
    inv02 ix36819 (.Y (nx36820), .A (nx37014)) ;
    inv02 ix36821 (.Y (nx36822), .A (nx37014)) ;
    inv02 ix36823 (.Y (nx36824), .A (nx37014)) ;
    inv02 ix36825 (.Y (nx36826), .A (nx37014)) ;
    inv02 ix36827 (.Y (nx36828), .A (nx8874)) ;
    inv02 ix36829 (.Y (nx36830), .A (nx37016)) ;
    inv02 ix36831 (.Y (nx36832), .A (nx37016)) ;
    inv02 ix36833 (.Y (nx36834), .A (nx37016)) ;
    inv02 ix36835 (.Y (nx36836), .A (nx37016)) ;
    inv02 ix36837 (.Y (nx36838), .A (nx37016)) ;
    inv02 ix36839 (.Y (nx36840), .A (nx11648)) ;
    inv02 ix36841 (.Y (nx36842), .A (nx37018)) ;
    inv02 ix36843 (.Y (nx36844), .A (nx37018)) ;
    inv02 ix36845 (.Y (nx36846), .A (nx37018)) ;
    inv02 ix36847 (.Y (nx36848), .A (nx37018)) ;
    inv02 ix36849 (.Y (nx36850), .A (nx37018)) ;
    inv02 ix36851 (.Y (nx36852), .A (nx14422)) ;
    inv02 ix36853 (.Y (nx36854), .A (nx37020)) ;
    inv02 ix36855 (.Y (nx36856), .A (nx37020)) ;
    inv02 ix36857 (.Y (nx36858), .A (nx37020)) ;
    inv02 ix36859 (.Y (nx36860), .A (nx37020)) ;
    inv02 ix36861 (.Y (nx36862), .A (nx37020)) ;
    inv02 ix36863 (.Y (nx36864), .A (nx17196)) ;
    inv02 ix36865 (.Y (nx36866), .A (nx37022)) ;
    inv02 ix36867 (.Y (nx36868), .A (nx37022)) ;
    inv02 ix36869 (.Y (nx36870), .A (nx37022)) ;
    inv02 ix36871 (.Y (nx36872), .A (nx37022)) ;
    inv02 ix36873 (.Y (nx36874), .A (nx37022)) ;
    inv02 ix36875 (.Y (nx36876), .A (nx19970)) ;
    inv02 ix36877 (.Y (nx36878), .A (nx37024)) ;
    inv02 ix36879 (.Y (nx36880), .A (nx37024)) ;
    inv02 ix36881 (.Y (nx36882), .A (nx37024)) ;
    inv02 ix36883 (.Y (nx36884), .A (nx37024)) ;
    inv02 ix36885 (.Y (nx36886), .A (nx37024)) ;
    inv02 ix36887 (.Y (nx36888), .A (nx22744)) ;
    inv02 ix36889 (.Y (nx36890), .A (nx37026)) ;
    inv02 ix36891 (.Y (nx36892), .A (nx37026)) ;
    inv02 ix36893 (.Y (nx36894), .A (nx37026)) ;
    inv02 ix36895 (.Y (nx36896), .A (nx37026)) ;
    inv02 ix36897 (.Y (nx36898), .A (nx37026)) ;
    inv04 ix36911 (.Y (nx36912), .A (nx37422)) ;
    inv02 ix36915 (.Y (nx36916), .A (nx23298)) ;
    inv02 ix36917 (.Y (nx36918), .A (nx23298)) ;
    inv02 ix36919 (.Y (nx36920), .A (nx23298)) ;
    inv02 ix36921 (.Y (nx36922), .A (nx36804)) ;
    inv02 ix36923 (.Y (nx36924), .A (nx23290)) ;
    inv02 ix36925 (.Y (nx36926), .A (nx23290)) ;
    inv02 ix36927 (.Y (nx36928), .A (nx23290)) ;
    inv02 ix36929 (.Y (nx36930), .A (nx23279)) ;
    inv02 ix36931 (.Y (nx36932), .A (nx23279)) ;
    inv02 ix36933 (.Y (nx36934), .A (nx23279)) ;
    inv02 ix36935 (.Y (nx36936), .A (nx23267)) ;
    inv02 ix36937 (.Y (nx36938), .A (nx23267)) ;
    inv02 ix36939 (.Y (nx36940), .A (nx23267)) ;
    inv02 ix36941 (.Y (nx36942), .A (nx36208)) ;
    inv02 ix36943 (.Y (nx36944), .A (nx36208)) ;
    inv02 ix36945 (.Y (nx36946), .A (nx36208)) ;
    inv02 ix36947 (.Y (nx36948), .A (nx36248)) ;
    inv02 ix36949 (.Y (nx36950), .A (nx36248)) ;
    inv02 ix36951 (.Y (nx36952), .A (nx36248)) ;
    inv02 ix36953 (.Y (nx36954), .A (nx36168)) ;
    inv02 ix36955 (.Y (nx36956), .A (nx36168)) ;
    inv02 ix36957 (.Y (nx36958), .A (nx36168)) ;
    inv02 ix36959 (.Y (nx36960), .A (nx36128)) ;
    inv02 ix36961 (.Y (nx36962), .A (nx36128)) ;
    inv02 ix36963 (.Y (nx36964), .A (nx36128)) ;
    inv02 ix36965 (.Y (nx36966), .A (nx36048)) ;
    inv02 ix36967 (.Y (nx36968), .A (nx36048)) ;
    inv02 ix36969 (.Y (nx36970), .A (nx36048)) ;
    inv02 ix36971 (.Y (nx36972), .A (nx36088)) ;
    inv02 ix36973 (.Y (nx36974), .A (nx36088)) ;
    inv02 ix36975 (.Y (nx36976), .A (nx36088)) ;
    inv02 ix36977 (.Y (nx36978), .A (nx36008)) ;
    inv02 ix36979 (.Y (nx36980), .A (nx36008)) ;
    inv02 ix36981 (.Y (nx36982), .A (nx36008)) ;
    inv02 ix36983 (.Y (nx36984), .A (nx35968)) ;
    inv02 ix36985 (.Y (nx36986), .A (nx35968)) ;
    inv02 ix36987 (.Y (nx36988), .A (nx35968)) ;
    inv02 ix36989 (.Y (nx36990), .A (nx35928)) ;
    inv02 ix36991 (.Y (nx36992), .A (nx35928)) ;
    inv02 ix36993 (.Y (nx36994), .A (nx35928)) ;
    inv02 ix36995 (.Y (nx36996), .A (nx35888)) ;
    inv02 ix36997 (.Y (nx36998), .A (nx35888)) ;
    inv02 ix36999 (.Y (nx37000), .A (nx35888)) ;
    inv02 ix37001 (.Y (nx37002), .A (nx35848)) ;
    inv02 ix37003 (.Y (nx37004), .A (nx35848)) ;
    inv02 ix37005 (.Y (nx37006), .A (nx35848)) ;
    inv02 ix37007 (.Y (nx37008), .A (nx35808)) ;
    inv02 ix37009 (.Y (nx37010), .A (nx35808)) ;
    inv02 ix37011 (.Y (nx37012), .A (nx35808)) ;
    inv02 ix37013 (.Y (nx37014), .A (nx36816)) ;
    inv02 ix37015 (.Y (nx37016), .A (nx36828)) ;
    inv02 ix37017 (.Y (nx37018), .A (nx36840)) ;
    inv02 ix37019 (.Y (nx37020), .A (nx36852)) ;
    inv02 ix37021 (.Y (nx37022), .A (nx36864)) ;
    inv02 ix37023 (.Y (nx37024), .A (nx36876)) ;
    inv02 ix37025 (.Y (nx37026), .A (nx36888)) ;
    inv04 ix37027 (.Y (nx37028), .A (camera_module_write_from_DMA)) ;
    inv02 ix37029 (.Y (nx37030), .A (nx1490)) ;
    inv02 ix37031 (.Y (nx37032), .A (nx1472)) ;
    inv02 ix37033 (.Y (nx37034), .A (nx1452)) ;
    inv02 ix37035 (.Y (nx37036), .A (nx1434)) ;
    inv02 ix37037 (.Y (nx37038), .A (nx1410)) ;
    inv02 ix37039 (.Y (nx37040), .A (nx1392)) ;
    inv02 ix37041 (.Y (nx37042), .A (nx1354)) ;
    inv02 ix37043 (.Y (nx37044), .A (nx1372)) ;
    inv02 ix37045 (.Y (nx37046), .A (nx1326)) ;
    inv02 ix37047 (.Y (nx37048), .A (nx1308)) ;
    inv02 ix37049 (.Y (nx37050), .A (nx1270)) ;
    inv02 ix37051 (.Y (nx37052), .A (nx1288)) ;
    mux21 ix27167 (.Y (nx27166), .A0 (nx35670), .A1 (motor_direction[0]), .S0 (
          nx37146)) ;
    and02 ix22580 (.Y (nx22579), .A0 (nx22585), .A1 (nx22943)) ;
    or03 ix22588 (.Y (nx22587), .A0 (rst), .A1 (nx22595), .A2 (nx35698)) ;
    mux21_ni ix1044 (.Y (nx1043), .A0 (camera_module_algo_module_pixel_enable), 
             .A1 (nx308), .S0 (nx879)) ;
    mux21_ni ix22524 (.Y (nx22523), .A0 (
             camera_module_algo_module_modCU_current_state_1), .A1 (nx27106), .S0 (
             nx879)) ;
    nor02ii ix27107 (.Y (nx27106), .A0 (rst), .A1 (nx37416)) ;
    nand04 ix22620 (.Y (nx879), .A0 (nx22565), .A1 (nx37058), .A2 (nx34018), .A3 (
           nx37060)) ;
    inv01 ix37057 (.Y (nx37058), .A (
          camera_module_algo_module_modCU_current_state_14)) ;
    inv01 ix37059 (.Y (nx37060), .A (nx27132)) ;
    xnor2 ix22632 (.Y (nx22631), .A0 (nx33810), .A1 (
          camera_module_algo_module_prev_cont_value_15)) ;
    mux21_ni ix22274 (.Y (nx22273), .A0 (
             camera_module_algo_module_current_cont_value_15), .A1 (nx26566), .S0 (
             nx37306)) ;
    mux21_ni ix26567 (.Y (nx26566), .A0 (
             camera_module_algo_module_Addout_value_15), .A1 (zero), .S0 (
             nx37074)) ;
    mux21_ni ix22264 (.Y (nx22263), .A0 (nx26552), .A1 (
             camera_module_algo_module_Addout_value_15), .S0 (nx37118)) ;
    mux21_ni ix26553 (.Y (nx26552), .A0 (zero), .A1 (nx26544), .S0 (nx37146)) ;
    mux21 ix22214 (.Y (nx22213), .A0 (nx22653), .A1 (nx22651), .S0 (nx37130)) ;
    oai21 ix22658 (.Y (nx25432), .A0 (nx33961), .A1 (nx37062), .B0 (nx22679)) ;
    inv01 ix37061 (.Y (nx37062), .A (nx22669)) ;
    and02 ix22666 (.Y (nx22665), .A0 (nx37136), .A1 (nx22601)) ;
    mux21 ix22609 (.Y (nx22608), .A0 (nx35674), .A1 (nx22699), .S0 (nx37136)) ;
    mux21_ni ix277 (.Y (nx276), .A0 (zero), .A1 (nx268), .S0 (nx37124)) ;
    mux21_ni ix227 (.Y (nx226), .A0 (zero), .A1 (nx218), .S0 (nx37124)) ;
    or04 ix22767 (.Y (nx22766), .A0 (nx22719), .A1 (nx37106), .A2 (nx37098), .A3 (
         nx37156)) ;
    mux21_ni ix22774 (.Y (nx22773), .A0 (nx35670), .A1 (nx22775), .S0 (nx37124)
             ) ;
    xor2 ix22778 (.Y (nx22777), .A0 (nx37106), .A1 (zero)) ;
    and02 ix22780 (.Y (nx22779), .A0 (nx37124), .A1 (nx37172)) ;
    mux21 ix22788 (.Y (nx22787), .A0 (zero), .A1 (nx56), .S0 (nx37126)) ;
    xor2 ix22792 (.Y (nx22791), .A0 (nx37156), .A1 (zero)) ;
    nor03_2x ix49 (.Y (nx48), .A0 (nx37064), .A1 (rst), .A2 (nx22611)) ;
    inv01 ix37063 (.Y (nx37064), .A (
          camera_module_DMA_module_controlUnit_state_1)) ;
    mux21 ix22806 (.Y (nx22805), .A0 (zero), .A1 (nx80), .S0 (nx37126)) ;
    ao22 ix79 (.Y (nx78), .A0 (zero), .A1 (nx37412), .B0 (one), .B1 (nx37066)) ;
    inv01 ix37065 (.Y (nx37066), .A (nx22791)) ;
    xor2 ix22812 (.Y (nx22811), .A0 (nx37098), .A1 (zero)) ;
    xor2 ix22816 (.Y (nx22815), .A0 (nx22821), .A1 (zero)) ;
    mux21_ni ix22824 (.Y (nx22823), .A0 (nx35670), .A1 (nx22825), .S0 (nx37126)
             ) ;
    xor2 ix22832 (.Y (nx22831), .A0 (nx22835), .A1 (zero)) ;
    mux21_ni ix22838 (.Y (nx22837), .A0 (nx35672), .A1 (nx22839), .S0 (nx37126)
             ) ;
    mux21 ix22847 (.Y (nx22846), .A0 (zero), .A1 (nx130), .S0 (nx37126)) ;
    xor2 ix22850 (.Y (nx22849), .A0 (nx22719), .A1 (zero)) ;
    mux21 ix22852 (.Y (nx22851), .A0 (nx19958), .A1 (nx19930), .S0 (nx37106)) ;
    mux21_ni ix19931 (.Y (nx19930), .A0 (nx19926), .A1 (nx19914), .S0 (nx37098)
             ) ;
    mux21_ni ix19915 (.Y (nx19914), .A0 (nvm_data_118), .A1 (nvm_data_126), .S0 (
             nx37158)) ;
    mux21_ni ix19927 (.Y (nx19926), .A0 (nvm_data_102), .A1 (nvm_data_110), .S0 (
             nx37158)) ;
    mux21_ni ix19959 (.Y (nx19958), .A0 (nx19954), .A1 (nx19942), .S0 (nx37098)
             ) ;
    mux21_ni ix19943 (.Y (nx19942), .A0 (nvm_data_86), .A1 (nvm_data_94), .S0 (
             nx37158)) ;
    mux21_ni ix19955 (.Y (nx19954), .A0 (nvm_data_70), .A1 (nvm_data_78), .S0 (
             nx37158)) ;
    mux21_ni ix19905 (.Y (nx19904), .A0 (nx19872), .A1 (nx19898), .S0 (nx37106)
             ) ;
    mux21_ni ix19899 (.Y (nx19898), .A0 (nx19894), .A1 (nx19882), .S0 (nx37098)
             ) ;
    mux21_ni ix19883 (.Y (nx19882), .A0 (nvm_data_54), .A1 (nvm_data_62), .S0 (
             nx37158)) ;
    mux21_ni ix19895 (.Y (nx19894), .A0 (nvm_data_38), .A1 (nvm_data_46), .S0 (
             nx37158)) ;
    mux21 ix22888 (.Y (nx22887), .A0 (nvm_data_22), .A1 (nvm_data_30), .S0 (
          nx37158)) ;
    and03 ix5921 (.Y (nx5920), .A0 (nx37200), .A1 (nx37436), .A2 (nx37232)) ;
    mux21_ni ix1051 (.Y (nx1050), .A0 (camera_module_cache_address_from_DMA_6), 
             .A1 (nx1042), .S0 (nx37172)) ;
    mux21_ni ix1043 (.Y (nx1042), .A0 (nx1032), .A1 (nx1038), .S0 (nx686)) ;
    xnor2 ix22908 (.Y (nx22907), .A0 (nx23011), .A1 (nx35782)) ;
    mux21_ni ix529 (.Y (nx528), .A0 (nx520), .A1 (zero), .S0 (nx37370)) ;
    mux21_ni ix471 (.Y (nx470), .A0 (nx462), .A1 (zero), .S0 (nx37370)) ;
    xnor2 ix22932 (.Y (nx22931), .A0 (nx22935), .A1 (nx35782)) ;
    mux21_ni ix1084 (.Y (nx1083), .A0 (
             camera_module_algo_module_modCU_current_state_7), .A1 (nx348), .S0 (
             nx879)) ;
    nor02ii ix349 (.Y (nx348), .A0 (rst), .A1 (
            camera_module_algo_module_modCU_current_state_6)) ;
    xor2 ix22952 (.Y (nx22951), .A0 (camera_module_algo_module_address_value_2)
         , .A1 (nx35782)) ;
    nor02ii ix22954 (.Y (nx22953), .A0 (
            camera_module_algo_module_prev_cont_enable), .A1 (nx37138)) ;
    mux21_ni ix22504 (.Y (nx22503), .A0 (motor_move), .A1 (nx27084), .S0 (nx879)
             ) ;
    mux21_ni ix27069 (.Y (nx27068), .A0 (zero), .A1 (one), .S0 (nx37138)) ;
    and02 ix22974 (.Y (nx22973), .A0 (nx37406), .A1 (nx22979)) ;
    or03 ix22982 (.Y (nx22981), .A0 (rst), .A1 (nx22987), .A2 (nx35698)) ;
    or03 ix22990 (.Y (nx22989), .A0 (rst), .A1 (nx22993), .A2 (nx35698)) ;
    xnor2 ix22998 (.Y (nx22997), .A0 (nx23005), .A1 (nx35782)) ;
    xor2 ix23007 (.Y (nx23006), .A0 (camera_module_algo_module_address_value_4)
         , .A1 (nx35782)) ;
    xor2 ix23027 (.Y (nx23026), .A0 (nx23021), .A1 (one)) ;
    xor2 ix23034 (.Y (nx23033), .A0 (camera_module_algo_module_address_value_6)
         , .A1 (nx35784)) ;
    mux21_ni ix577 (.Y (nx576), .A0 (nx568), .A1 (zero), .S0 (nx37370)) ;
    mux21_ni ix1033 (.Y (nx1032), .A0 (camera_module_algo_module_address_value_6
             ), .A1 (nx568), .S0 (nx37082)) ;
    nand02 ix23044 (.Y (nx688), .A0 (nx22597), .A1 (nx22943)) ;
    nand02_2x ix23047 (.Y (nx686), .A0 (nx22585), .A1 (nx22987)) ;
    mux21_ni ix1025 (.Y (nx1024), .A0 (camera_module_cache_address_from_DMA_7), 
             .A1 (nx1016), .S0 (nx37172)) ;
    mux21_ni ix23052 (.Y (nx23051), .A0 (nx23067), .A1 (nx23053), .S0 (nx37082)
             ) ;
    xnor2 ix23060 (.Y (nx23059), .A0 (nx23067), .A1 (nx35784)) ;
    mux21_ni ix981 (.Y (nx980), .A0 (camera_module_cache_address_from_DMA_4), .A1 (
             nx972), .S0 (nx37172)) ;
    mux21_ni ix973 (.Y (nx972), .A0 (nx962), .A1 (nx968), .S0 (nx686)) ;
    mux21_ni ix963 (.Y (nx962), .A0 (camera_module_algo_module_address_value_4)
             , .A1 (nx520), .S0 (nx37082)) ;
    mux21_ni ix955 (.Y (nx954), .A0 (camera_module_cache_address_from_DMA_5), .A1 (
             nx946), .S0 (nx37172)) ;
    mux21_ni ix23085 (.Y (nx23084), .A0 (nx23011), .A1 (nx22912), .S0 (nx37082)
             ) ;
    mux21_ni ix907 (.Y (nx906), .A0 (nx34112), .A1 (nx898), .S0 (nx37174)) ;
    mux21_ni ix899 (.Y (nx898), .A0 (nx888), .A1 (nx894), .S0 (nx686)) ;
    mux21_ni ix889 (.Y (nx888), .A0 (camera_module_algo_module_address_value_2)
             , .A1 (nx462), .S0 (nx37084)) ;
    mux21_ni ix881 (.Y (nx880), .A0 (nx34072), .A1 (nx872), .S0 (nx37174)) ;
    mux21_ni ix23101 (.Y (nx23100), .A0 (nx23005), .A1 (nx23003), .S0 (nx37084)
             ) ;
    mux21_ni ix837 (.Y (nx836), .A0 (nx34080), .A1 (nx828), .S0 (nx37174)) ;
    mux21_ni ix23112 (.Y (nx23111), .A0 (nx23021), .A1 (nx23026), .S0 (nx37084)
             ) ;
    xor2 ix23114 (.Y (nx23113), .A0 (nx23021), .A1 (zero)) ;
    mux21_ni ix811 (.Y (nx810), .A0 (nx34100), .A1 (nx802), .S0 (nx37174)) ;
    mux21_ni ix23118 (.Y (nx23117), .A0 (nx22935), .A1 (nx22575), .S0 (nx37084)
             ) ;
    and03 ix5905 (.Y (nx5904), .A0 (nx37202), .A1 (nx37436), .A2 (nx37232)) ;
    nor02ii ix23131 (.Y (nx23130), .A0 (nx954), .A1 (nx980)) ;
    and03 ix5887 (.Y (nx5886), .A0 (nx37204), .A1 (nx37436), .A2 (nx37232)) ;
    nor02ii ix23146 (.Y (nx23145), .A0 (nx980), .A1 (nx954)) ;
    and03 ix5871 (.Y (nx5870), .A0 (nx37206), .A1 (nx37436), .A2 (nx37232)) ;
    and03 ix5851 (.Y (nx5850), .A0 (nx37208), .A1 (nx37436), .A2 (nx37232)) ;
    nor02ii ix23173 (.Y (nx23172), .A0 (nx1024), .A1 (nx1050)) ;
    and03 ix5835 (.Y (nx5834), .A0 (nx37210), .A1 (nx37436), .A2 (nx37232)) ;
    and03 ix5801 (.Y (nx5800), .A0 (nx37212), .A1 (nx37312), .A2 (nx37234)) ;
    and03 ix5817 (.Y (nx5816), .A0 (nx37214), .A1 (nx37312), .A2 (nx37234)) ;
    and03 ix5779 (.Y (nx5778), .A0 (nx37216), .A1 (nx37312), .A2 (nx37234)) ;
    nor02ii ix23219 (.Y (nx23218), .A0 (nx1050), .A1 (nx1024)) ;
    and03 ix5763 (.Y (nx5762), .A0 (nx37218), .A1 (nx37312), .A2 (nx37234)) ;
    and03 ix5729 (.Y (nx5728), .A0 (nx37220), .A1 (nx37312), .A2 (nx37234)) ;
    and03 ix5745 (.Y (nx5744), .A0 (nx37222), .A1 (nx37312), .A2 (nx37234)) ;
    and03 ix5709 (.Y (nx5708), .A0 (nx37224), .A1 (nx37312), .A2 (nx37234)) ;
    nor02ii ix23268 (.Y (nx23267), .A0 (nx1056), .A1 (nx23073)) ;
    and03 ix5693 (.Y (nx5692), .A0 (nx37226), .A1 (nx37314), .A2 (nx36450)) ;
    nor02ii ix23280 (.Y (nx23279), .A0 (nx1056), .A1 (nx23130)) ;
    and03 ix5675 (.Y (nx5674), .A0 (nx37228), .A1 (nx37314), .A2 (nx36450)) ;
    nor02ii ix23291 (.Y (nx23290), .A0 (nx1056), .A1 (nx23145)) ;
    and03 ix5659 (.Y (nx5658), .A0 (nx37230), .A1 (nx37314), .A2 (nx36450)) ;
    and03 ix5629 (.Y (nx5628), .A0 (nx37236), .A1 (nx37314), .A2 (nx35844)) ;
    nor02ii ix23315 (.Y (nx23314), .A0 (nx810), .A1 (nx836)) ;
    and03 ix5613 (.Y (nx5612), .A0 (nx35884), .A1 (nx37314), .A2 (nx37236)) ;
    and03 ix5595 (.Y (nx5594), .A0 (nx35924), .A1 (nx37314), .A2 (nx37236)) ;
    and03 ix5579 (.Y (nx5578), .A0 (nx35964), .A1 (nx37314), .A2 (nx37236)) ;
    and03 ix5559 (.Y (nx5558), .A0 (nx36004), .A1 (nx37316), .A2 (nx37236)) ;
    and03 ix5543 (.Y (nx5542), .A0 (nx36044), .A1 (nx37316), .A2 (nx37236)) ;
    and03 ix5509 (.Y (nx5508), .A0 (nx36084), .A1 (nx37316), .A2 (nx37238)) ;
    and03 ix5525 (.Y (nx5524), .A0 (nx36124), .A1 (nx37316), .A2 (nx37238)) ;
    and03 ix5487 (.Y (nx5486), .A0 (nx36164), .A1 (nx37316), .A2 (nx37238)) ;
    and03 ix5471 (.Y (nx5470), .A0 (nx36204), .A1 (nx37316), .A2 (nx37238)) ;
    and03 ix5437 (.Y (nx5436), .A0 (nx36244), .A1 (nx37316), .A2 (nx37238)) ;
    and03 ix5453 (.Y (nx5452), .A0 (nx36284), .A1 (nx37318), .A2 (nx37238)) ;
    and03 ix5417 (.Y (nx5416), .A0 (nx36324), .A1 (nx37318), .A2 (nx37238)) ;
    and03 ix5401 (.Y (nx5400), .A0 (nx36364), .A1 (nx37318), .A2 (nx36454)) ;
    and03 ix5383 (.Y (nx5382), .A0 (nx36404), .A1 (nx37318), .A2 (nx36454)) ;
    and03 ix5367 (.Y (nx5366), .A0 (nx36444), .A1 (nx37318), .A2 (nx36454)) ;
    and03 ix5335 (.Y (nx5334), .A0 (nx37240), .A1 (nx37318), .A2 (nx35844)) ;
    nor02ii ix23424 (.Y (nx23423), .A0 (nx836), .A1 (nx810)) ;
    and03 ix5319 (.Y (nx5318), .A0 (nx35884), .A1 (nx37318), .A2 (nx37240)) ;
    and03 ix5301 (.Y (nx5300), .A0 (nx35924), .A1 (nx37320), .A2 (nx37240)) ;
    and03 ix5285 (.Y (nx5284), .A0 (nx35964), .A1 (nx37320), .A2 (nx37240)) ;
    and03 ix5265 (.Y (nx5264), .A0 (nx36004), .A1 (nx37320), .A2 (nx37240)) ;
    and03 ix5249 (.Y (nx5248), .A0 (nx36044), .A1 (nx37320), .A2 (nx37240)) ;
    and03 ix5215 (.Y (nx5214), .A0 (nx36084), .A1 (nx37320), .A2 (nx37242)) ;
    and03 ix5231 (.Y (nx5230), .A0 (nx36124), .A1 (nx37320), .A2 (nx37242)) ;
    and03 ix5193 (.Y (nx5192), .A0 (nx36164), .A1 (nx37320), .A2 (nx37242)) ;
    and03 ix5177 (.Y (nx5176), .A0 (nx36204), .A1 (nx37322), .A2 (nx37242)) ;
    and03 ix5143 (.Y (nx5142), .A0 (nx36244), .A1 (nx37322), .A2 (nx37242)) ;
    and03 ix5159 (.Y (nx5158), .A0 (nx36284), .A1 (nx37322), .A2 (nx37242)) ;
    and03 ix5123 (.Y (nx5122), .A0 (nx36324), .A1 (nx37322), .A2 (nx37242)) ;
    and03 ix5107 (.Y (nx5106), .A0 (nx36364), .A1 (nx37322), .A2 (nx36458)) ;
    and03 ix5089 (.Y (nx5088), .A0 (nx36404), .A1 (nx37322), .A2 (nx36458)) ;
    and03 ix5073 (.Y (nx5072), .A0 (nx36444), .A1 (nx37322), .A2 (nx36458)) ;
    and03 ix5043 (.Y (nx5042), .A0 (nx37244), .A1 (nx37324), .A2 (nx35844)) ;
    and03 ix5027 (.Y (nx5026), .A0 (nx35884), .A1 (nx37324), .A2 (nx37244)) ;
    and03 ix5009 (.Y (nx5008), .A0 (nx35924), .A1 (nx37324), .A2 (nx37244)) ;
    and03 ix4993 (.Y (nx4992), .A0 (nx35964), .A1 (nx37324), .A2 (nx37244)) ;
    and03 ix4973 (.Y (nx4972), .A0 (nx36004), .A1 (nx37324), .A2 (nx37244)) ;
    and03 ix4957 (.Y (nx4956), .A0 (nx36044), .A1 (nx37324), .A2 (nx37244)) ;
    and03 ix4923 (.Y (nx4922), .A0 (nx36084), .A1 (nx37324), .A2 (nx37246)) ;
    and03 ix4939 (.Y (nx4938), .A0 (nx36124), .A1 (nx37326), .A2 (nx37246)) ;
    and03 ix4901 (.Y (nx4900), .A0 (nx36164), .A1 (nx37326), .A2 (nx37246)) ;
    and03 ix4885 (.Y (nx4884), .A0 (nx36204), .A1 (nx37326), .A2 (nx37246)) ;
    and03 ix4851 (.Y (nx4850), .A0 (nx36244), .A1 (nx37326), .A2 (nx37246)) ;
    and03 ix4867 (.Y (nx4866), .A0 (nx36284), .A1 (nx37326), .A2 (nx37246)) ;
    and03 ix4831 (.Y (nx4830), .A0 (nx36324), .A1 (nx37326), .A2 (nx37246)) ;
    and03 ix4815 (.Y (nx4814), .A0 (nx36364), .A1 (nx37326), .A2 (nx36462)) ;
    and03 ix4797 (.Y (nx4796), .A0 (nx36404), .A1 (nx37328), .A2 (nx36462)) ;
    and03 ix4781 (.Y (nx4780), .A0 (nx36444), .A1 (nx37328), .A2 (nx36462)) ;
    and03 ix4745 (.Y (nx4744), .A0 (nx37248), .A1 (nx37328), .A2 (nx35844)) ;
    nor02ii ix23640 (.Y (nx23639), .A0 (nx880), .A1 (nx906)) ;
    and03 ix4729 (.Y (nx4728), .A0 (nx35884), .A1 (nx37328), .A2 (nx37248)) ;
    and03 ix4711 (.Y (nx4710), .A0 (nx35924), .A1 (nx37328), .A2 (nx37248)) ;
    and03 ix4695 (.Y (nx4694), .A0 (nx35964), .A1 (nx37328), .A2 (nx37248)) ;
    and03 ix4675 (.Y (nx4674), .A0 (nx36004), .A1 (nx37328), .A2 (nx37248)) ;
    and03 ix4659 (.Y (nx4658), .A0 (nx36044), .A1 (nx37330), .A2 (nx37248)) ;
    and03 ix4625 (.Y (nx4624), .A0 (nx36084), .A1 (nx37330), .A2 (nx37250)) ;
    and03 ix4641 (.Y (nx4640), .A0 (nx36124), .A1 (nx37330), .A2 (nx37250)) ;
    and03 ix4603 (.Y (nx4602), .A0 (nx36164), .A1 (nx37330), .A2 (nx37250)) ;
    and03 ix4587 (.Y (nx4586), .A0 (nx36204), .A1 (nx37330), .A2 (nx37250)) ;
    and03 ix4553 (.Y (nx4552), .A0 (nx36244), .A1 (nx37330), .A2 (nx37250)) ;
    and03 ix4569 (.Y (nx4568), .A0 (nx36284), .A1 (nx37330), .A2 (nx37250)) ;
    and03 ix4533 (.Y (nx4532), .A0 (nx36324), .A1 (nx37332), .A2 (nx37250)) ;
    and03 ix4517 (.Y (nx4516), .A0 (nx36364), .A1 (nx37332), .A2 (nx36466)) ;
    and03 ix4499 (.Y (nx4498), .A0 (nx36404), .A1 (nx37332), .A2 (nx36466)) ;
    and03 ix4483 (.Y (nx4482), .A0 (nx36444), .A1 (nx37332), .A2 (nx36466)) ;
    and03 ix4453 (.Y (nx4452), .A0 (nx37252), .A1 (nx37332), .A2 (nx35844)) ;
    and03 ix4437 (.Y (nx4436), .A0 (nx35884), .A1 (nx37332), .A2 (nx37252)) ;
    and03 ix4419 (.Y (nx4418), .A0 (nx35924), .A1 (nx37332), .A2 (nx37252)) ;
    and03 ix4403 (.Y (nx4402), .A0 (nx35964), .A1 (nx37334), .A2 (nx37252)) ;
    and03 ix4383 (.Y (nx4382), .A0 (nx36004), .A1 (nx37334), .A2 (nx37252)) ;
    and03 ix4367 (.Y (nx4366), .A0 (nx36044), .A1 (nx37334), .A2 (nx37252)) ;
    and03 ix4333 (.Y (nx4332), .A0 (nx36084), .A1 (nx37334), .A2 (nx37254)) ;
    and03 ix4349 (.Y (nx4348), .A0 (nx36124), .A1 (nx37334), .A2 (nx37254)) ;
    and03 ix4311 (.Y (nx4310), .A0 (nx36164), .A1 (nx37334), .A2 (nx37254)) ;
    and03 ix4295 (.Y (nx4294), .A0 (nx36204), .A1 (nx37334), .A2 (nx37254)) ;
    and03 ix4261 (.Y (nx4260), .A0 (nx36244), .A1 (nx37336), .A2 (nx37254)) ;
    and03 ix4277 (.Y (nx4276), .A0 (nx36284), .A1 (nx37336), .A2 (nx37254)) ;
    and03 ix4241 (.Y (nx4240), .A0 (nx36324), .A1 (nx37336), .A2 (nx37254)) ;
    and03 ix4225 (.Y (nx4224), .A0 (nx36364), .A1 (nx37336), .A2 (nx36470)) ;
    and03 ix4207 (.Y (nx4206), .A0 (nx36404), .A1 (nx37336), .A2 (nx36470)) ;
    and03 ix4191 (.Y (nx4190), .A0 (nx36444), .A1 (nx37336), .A2 (nx36470)) ;
    and03 ix4159 (.Y (nx4158), .A0 (nx37256), .A1 (nx37336), .A2 (nx35846)) ;
    and03 ix4143 (.Y (nx4142), .A0 (nx35884), .A1 (nx37338), .A2 (nx37256)) ;
    and03 ix4125 (.Y (nx4124), .A0 (nx35924), .A1 (nx37338), .A2 (nx37256)) ;
    and03 ix4109 (.Y (nx4108), .A0 (nx35964), .A1 (nx37338), .A2 (nx37256)) ;
    and03 ix4089 (.Y (nx4088), .A0 (nx36004), .A1 (nx37338), .A2 (nx37256)) ;
    and03 ix4073 (.Y (nx4072), .A0 (nx36044), .A1 (nx37338), .A2 (nx37256)) ;
    and03 ix4039 (.Y (nx4038), .A0 (nx36084), .A1 (nx37338), .A2 (nx37258)) ;
    and03 ix4055 (.Y (nx4054), .A0 (nx36124), .A1 (nx37338), .A2 (nx37258)) ;
    and03 ix4017 (.Y (nx4016), .A0 (nx36164), .A1 (nx37340), .A2 (nx37258)) ;
    and03 ix4001 (.Y (nx4000), .A0 (nx36204), .A1 (nx37340), .A2 (nx37258)) ;
    and03 ix3967 (.Y (nx3966), .A0 (nx36244), .A1 (nx37340), .A2 (nx37258)) ;
    and03 ix3983 (.Y (nx3982), .A0 (nx36284), .A1 (nx37340), .A2 (nx37258)) ;
    and03 ix3947 (.Y (nx3946), .A0 (nx36324), .A1 (nx37340), .A2 (nx37258)) ;
    and03 ix3931 (.Y (nx3930), .A0 (nx36364), .A1 (nx37340), .A2 (nx36474)) ;
    and03 ix3913 (.Y (nx3912), .A0 (nx36404), .A1 (nx37340), .A2 (nx36474)) ;
    and03 ix3897 (.Y (nx3896), .A0 (nx36444), .A1 (nx37342), .A2 (nx36474)) ;
    and03 ix3867 (.Y (nx3866), .A0 (nx37260), .A1 (nx37342), .A2 (nx35846)) ;
    and03 ix3851 (.Y (nx3850), .A0 (nx35886), .A1 (nx37342), .A2 (nx37260)) ;
    and03 ix3833 (.Y (nx3832), .A0 (nx35926), .A1 (nx37342), .A2 (nx37260)) ;
    and03 ix3817 (.Y (nx3816), .A0 (nx35966), .A1 (nx37342), .A2 (nx37260)) ;
    and03 ix3797 (.Y (nx3796), .A0 (nx36006), .A1 (nx37342), .A2 (nx37260)) ;
    and03 ix3781 (.Y (nx3780), .A0 (nx36046), .A1 (nx37342), .A2 (nx37260)) ;
    and03 ix3747 (.Y (nx3746), .A0 (nx36086), .A1 (nx37344), .A2 (nx37262)) ;
    and03 ix3763 (.Y (nx3762), .A0 (nx36126), .A1 (nx37344), .A2 (nx37262)) ;
    and03 ix3725 (.Y (nx3724), .A0 (nx36166), .A1 (nx37344), .A2 (nx37262)) ;
    and03 ix3709 (.Y (nx3708), .A0 (nx36206), .A1 (nx37344), .A2 (nx37262)) ;
    and03 ix3675 (.Y (nx3674), .A0 (nx36246), .A1 (nx37344), .A2 (nx37262)) ;
    and03 ix3691 (.Y (nx3690), .A0 (nx36286), .A1 (nx37344), .A2 (nx37262)) ;
    and03 ix3655 (.Y (nx3654), .A0 (nx36326), .A1 (nx37344), .A2 (nx37262)) ;
    and03 ix3639 (.Y (nx3638), .A0 (nx36366), .A1 (nx37346), .A2 (nx36478)) ;
    and03 ix3621 (.Y (nx3620), .A0 (nx36406), .A1 (nx37346), .A2 (nx36478)) ;
    and03 ix3605 (.Y (nx3604), .A0 (nx36446), .A1 (nx37346), .A2 (nx36478)) ;
    and03 ix3565 (.Y (nx3564), .A0 (nx37264), .A1 (nx37346), .A2 (nx35846)) ;
    nor02ii ix24054 (.Y (nx24053), .A0 (nx906), .A1 (nx880)) ;
    and03 ix3549 (.Y (nx3548), .A0 (nx35886), .A1 (nx37346), .A2 (nx37264)) ;
    and03 ix3531 (.Y (nx3530), .A0 (nx35926), .A1 (nx37346), .A2 (nx37264)) ;
    and03 ix3515 (.Y (nx3514), .A0 (nx35966), .A1 (nx37346), .A2 (nx37264)) ;
    and03 ix3495 (.Y (nx3494), .A0 (nx36006), .A1 (nx37348), .A2 (nx37264)) ;
    and03 ix3479 (.Y (nx3478), .A0 (nx36046), .A1 (nx37348), .A2 (nx37264)) ;
    and03 ix3445 (.Y (nx3444), .A0 (nx36086), .A1 (nx37348), .A2 (nx37266)) ;
    and03 ix3461 (.Y (nx3460), .A0 (nx36126), .A1 (nx37348), .A2 (nx37266)) ;
    and03 ix3423 (.Y (nx3422), .A0 (nx36166), .A1 (nx37348), .A2 (nx37266)) ;
    and03 ix3407 (.Y (nx3406), .A0 (nx36206), .A1 (nx37348), .A2 (nx37266)) ;
    and03 ix3373 (.Y (nx3372), .A0 (nx36246), .A1 (nx37348), .A2 (nx37266)) ;
    and03 ix3389 (.Y (nx3388), .A0 (nx36286), .A1 (nx37350), .A2 (nx37266)) ;
    and03 ix3353 (.Y (nx3352), .A0 (nx36326), .A1 (nx37350), .A2 (nx37266)) ;
    and03 ix3337 (.Y (nx3336), .A0 (nx36366), .A1 (nx37350), .A2 (nx36482)) ;
    and03 ix3319 (.Y (nx3318), .A0 (nx36406), .A1 (nx37350), .A2 (nx36482)) ;
    and03 ix3303 (.Y (nx3302), .A0 (nx36446), .A1 (nx37350), .A2 (nx36482)) ;
    and03 ix3273 (.Y (nx3272), .A0 (nx37268), .A1 (nx37350), .A2 (nx35846)) ;
    and03 ix3257 (.Y (nx3256), .A0 (nx35886), .A1 (nx37350), .A2 (nx37268)) ;
    and03 ix3239 (.Y (nx3238), .A0 (nx35926), .A1 (nx37352), .A2 (nx37268)) ;
    and03 ix3223 (.Y (nx3222), .A0 (nx35966), .A1 (nx37352), .A2 (nx37268)) ;
    and03 ix3203 (.Y (nx3202), .A0 (nx36006), .A1 (nx37352), .A2 (nx37268)) ;
    and03 ix3187 (.Y (nx3186), .A0 (nx36046), .A1 (nx37352), .A2 (nx37268)) ;
    and03 ix3153 (.Y (nx3152), .A0 (nx36086), .A1 (nx37352), .A2 (nx37270)) ;
    and03 ix3169 (.Y (nx3168), .A0 (nx36126), .A1 (nx37352), .A2 (nx37270)) ;
    and03 ix3131 (.Y (nx3130), .A0 (nx36166), .A1 (nx37352), .A2 (nx37270)) ;
    and03 ix3115 (.Y (nx3114), .A0 (nx36206), .A1 (nx37354), .A2 (nx37270)) ;
    and03 ix3081 (.Y (nx3080), .A0 (nx36246), .A1 (nx37354), .A2 (nx37270)) ;
    and03 ix3097 (.Y (nx3096), .A0 (nx36286), .A1 (nx37354), .A2 (nx37270)) ;
    and03 ix3061 (.Y (nx3060), .A0 (nx36326), .A1 (nx37354), .A2 (nx37270)) ;
    and03 ix3045 (.Y (nx3044), .A0 (nx36366), .A1 (nx37354), .A2 (nx36486)) ;
    and03 ix3027 (.Y (nx3026), .A0 (nx36406), .A1 (nx37356), .A2 (nx36486)) ;
    and03 ix3011 (.Y (nx3010), .A0 (nx36446), .A1 (nx37356), .A2 (nx36486)) ;
    and03 ix2979 (.Y (nx2978), .A0 (nx37272), .A1 (nx37356), .A2 (nx35846)) ;
    and03 ix2963 (.Y (nx2962), .A0 (nx35886), .A1 (nx37356), .A2 (nx37272)) ;
    and03 ix2945 (.Y (nx2944), .A0 (nx35926), .A1 (nx37356), .A2 (nx37272)) ;
    and03 ix2929 (.Y (nx2928), .A0 (nx35966), .A1 (nx37356), .A2 (nx37272)) ;
    and03 ix2909 (.Y (nx2908), .A0 (nx36006), .A1 (nx37356), .A2 (nx37272)) ;
    and03 ix2893 (.Y (nx2892), .A0 (nx36046), .A1 (nx37358), .A2 (nx37272)) ;
    and03 ix2859 (.Y (nx2858), .A0 (nx36086), .A1 (nx37358), .A2 (nx37274)) ;
    and03 ix2875 (.Y (nx2874), .A0 (nx36126), .A1 (nx37358), .A2 (nx37274)) ;
    and03 ix2837 (.Y (nx2836), .A0 (nx36166), .A1 (nx37358), .A2 (nx37274)) ;
    and03 ix2821 (.Y (nx2820), .A0 (nx36206), .A1 (nx37358), .A2 (nx37274)) ;
    and03 ix2787 (.Y (nx2786), .A0 (nx36246), .A1 (nx37358), .A2 (nx37274)) ;
    and03 ix2803 (.Y (nx2802), .A0 (nx36286), .A1 (nx37358), .A2 (nx37274)) ;
    and03 ix2767 (.Y (nx2766), .A0 (nx36326), .A1 (nx37360), .A2 (nx37274)) ;
    and03 ix2751 (.Y (nx2750), .A0 (nx36366), .A1 (nx37360), .A2 (nx36490)) ;
    and03 ix2733 (.Y (nx2732), .A0 (nx36406), .A1 (nx37360), .A2 (nx36490)) ;
    and03 ix2717 (.Y (nx2716), .A0 (nx36446), .A1 (nx37360), .A2 (nx36490)) ;
    and03 ix2687 (.Y (nx2686), .A0 (nx37276), .A1 (nx37360), .A2 (nx35846)) ;
    and03 ix2671 (.Y (nx2670), .A0 (nx35886), .A1 (nx37360), .A2 (nx37276)) ;
    and03 ix2653 (.Y (nx2652), .A0 (nx35926), .A1 (nx37360), .A2 (nx37276)) ;
    and03 ix2637 (.Y (nx2636), .A0 (nx35966), .A1 (nx37362), .A2 (nx37276)) ;
    and03 ix2617 (.Y (nx2616), .A0 (nx36006), .A1 (nx37362), .A2 (nx37276)) ;
    and03 ix2601 (.Y (nx2600), .A0 (nx36046), .A1 (nx37362), .A2 (nx37276)) ;
    and03 ix2567 (.Y (nx2566), .A0 (nx36086), .A1 (nx37362), .A2 (nx37278)) ;
    and03 ix2583 (.Y (nx2582), .A0 (nx36126), .A1 (nx37362), .A2 (nx37278)) ;
    and03 ix2545 (.Y (nx2544), .A0 (nx36166), .A1 (nx37362), .A2 (nx37278)) ;
    and03 ix2529 (.Y (nx2528), .A0 (nx36206), .A1 (nx37362), .A2 (nx37278)) ;
    and03 ix2495 (.Y (nx2494), .A0 (nx36246), .A1 (nx37364), .A2 (nx37278)) ;
    and03 ix2511 (.Y (nx2510), .A0 (nx36286), .A1 (nx37364), .A2 (nx37278)) ;
    and03 ix2475 (.Y (nx2474), .A0 (nx36326), .A1 (nx37364), .A2 (nx37278)) ;
    and03 ix2459 (.Y (nx2458), .A0 (nx36366), .A1 (nx37364), .A2 (nx36494)) ;
    and03 ix2441 (.Y (nx2440), .A0 (nx36406), .A1 (nx37364), .A2 (nx36494)) ;
    and03 ix2425 (.Y (nx2424), .A0 (nx36446), .A1 (nx37364), .A2 (nx36494)) ;
    or03 ix24464 (.Y (nx24463), .A0 (nx37280), .A1 (nx37174), .A2 (nx37008)) ;
    nand02 ix24466 (.Y (nx36500), .A0 (nx37068), .A1 (nx23105)) ;
    inv01 ix37067 (.Y (nx37068), .A (nx912)) ;
    or03 ix24474 (.Y (nx24473), .A0 (nx37002), .A1 (nx37174), .A2 (nx37280)) ;
    or03 ix24482 (.Y (nx24481), .A0 (nx36996), .A1 (nx37174), .A2 (nx37280)) ;
    or03 ix24488 (.Y (nx24487), .A0 (nx36990), .A1 (nx37176), .A2 (nx37280)) ;
    or03 ix24496 (.Y (nx24495), .A0 (nx36984), .A1 (nx37176), .A2 (nx37280)) ;
    or03 ix24501 (.Y (nx24500), .A0 (nx36978), .A1 (nx37178), .A2 (nx37280)) ;
    or03 ix24509 (.Y (nx24508), .A0 (nx36966), .A1 (nx37178), .A2 (nx37282)) ;
    or03 ix24514 (.Y (nx24513), .A0 (nx36972), .A1 (nx37178), .A2 (nx37282)) ;
    or03 ix24522 (.Y (nx24521), .A0 (nx36960), .A1 (nx37178), .A2 (nx37282)) ;
    or03 ix24527 (.Y (nx24526), .A0 (nx36954), .A1 (nx37178), .A2 (nx37282)) ;
    or03 ix24536 (.Y (nx24535), .A0 (nx36942), .A1 (nx37178), .A2 (nx37282)) ;
    or03 ix24542 (.Y (nx24541), .A0 (nx36948), .A1 (nx37178), .A2 (nx37282)) ;
    or03 ix24549 (.Y (nx24548), .A0 (nx36936), .A1 (nx37180), .A2 (nx37282)) ;
    or03 ix24555 (.Y (nx24554), .A0 (nx36930), .A1 (nx37180), .A2 (nx37284)) ;
    or03 ix24564 (.Y (nx24563), .A0 (nx36924), .A1 (nx37180), .A2 (nx37284)) ;
    or03 ix24570 (.Y (nx24569), .A0 (nx36916), .A1 (nx37180), .A2 (nx37284)) ;
    or03 ix24582 (.Y (nx24581), .A0 (nx37286), .A1 (nx37180), .A2 (nx37008)) ;
    nand02 ix24584 (.Y (nx36574), .A0 (nx37068), .A1 (nx23314)) ;
    or03 ix24590 (.Y (nx24589), .A0 (nx37002), .A1 (nx37180), .A2 (nx37286)) ;
    or03 ix24598 (.Y (nx24597), .A0 (nx36996), .A1 (nx37180), .A2 (nx37286)) ;
    or03 ix24603 (.Y (nx24602), .A0 (nx36990), .A1 (nx37182), .A2 (nx37286)) ;
    or03 ix24611 (.Y (nx24610), .A0 (nx36984), .A1 (nx37182), .A2 (nx37286)) ;
    or03 ix24616 (.Y (nx24615), .A0 (nx36978), .A1 (nx37182), .A2 (nx37286)) ;
    or03 ix24625 (.Y (nx24624), .A0 (nx36966), .A1 (nx37182), .A2 (nx37288)) ;
    or03 ix24630 (.Y (nx24629), .A0 (nx36972), .A1 (nx37182), .A2 (nx37288)) ;
    or03 ix24638 (.Y (nx24637), .A0 (nx36960), .A1 (nx37182), .A2 (nx37288)) ;
    or03 ix24643 (.Y (nx24642), .A0 (nx36954), .A1 (nx37182), .A2 (nx37288)) ;
    or03 ix24651 (.Y (nx24650), .A0 (nx36942), .A1 (nx37184), .A2 (nx37288)) ;
    or03 ix24656 (.Y (nx24655), .A0 (nx36948), .A1 (nx37184), .A2 (nx37288)) ;
    or03 ix24664 (.Y (nx24663), .A0 (nx36936), .A1 (nx37184), .A2 (nx37288)) ;
    or03 ix24670 (.Y (nx24669), .A0 (nx36930), .A1 (nx37184), .A2 (nx37290)) ;
    or03 ix24678 (.Y (nx24677), .A0 (nx36924), .A1 (nx37184), .A2 (nx37290)) ;
    or03 ix24683 (.Y (nx24682), .A0 (nx36916), .A1 (nx37184), .A2 (nx37290)) ;
    or03 ix24694 (.Y (nx24693), .A0 (nx37292), .A1 (nx37184), .A2 (nx37008)) ;
    nand02 ix24696 (.Y (nx36648), .A0 (nx37068), .A1 (nx23423)) ;
    or03 ix24704 (.Y (nx24703), .A0 (nx37002), .A1 (nx37186), .A2 (nx37292)) ;
    or03 ix24713 (.Y (nx24712), .A0 (nx36996), .A1 (nx37186), .A2 (nx37292)) ;
    or03 ix24718 (.Y (nx24717), .A0 (nx36990), .A1 (nx37186), .A2 (nx37292)) ;
    or03 ix24726 (.Y (nx24725), .A0 (nx36984), .A1 (nx37186), .A2 (nx37292)) ;
    or03 ix24731 (.Y (nx24730), .A0 (nx36978), .A1 (nx37186), .A2 (nx37292)) ;
    or03 ix24739 (.Y (nx24738), .A0 (nx36966), .A1 (nx37186), .A2 (nx37294)) ;
    or03 ix24744 (.Y (nx24743), .A0 (nx36972), .A1 (nx37186), .A2 (nx37294)) ;
    or03 ix24752 (.Y (nx24751), .A0 (nx36960), .A1 (nx37188), .A2 (nx37294)) ;
    or03 ix24758 (.Y (nx24757), .A0 (nx36954), .A1 (nx37188), .A2 (nx37294)) ;
    or03 ix24766 (.Y (nx24765), .A0 (nx36942), .A1 (nx37188), .A2 (nx37294)) ;
    or03 ix24771 (.Y (nx24770), .A0 (nx36948), .A1 (nx37188), .A2 (nx37294)) ;
    or03 ix24779 (.Y (nx24778), .A0 (nx36936), .A1 (nx37188), .A2 (nx37294)) ;
    or03 ix24786 (.Y (nx24785), .A0 (nx36930), .A1 (nx37188), .A2 (nx37296)) ;
    or03 ix24793 (.Y (nx24792), .A0 (nx36924), .A1 (nx37188), .A2 (nx37296)) ;
    or03 ix24799 (.Y (nx24798), .A0 (nx36916), .A1 (nx37190), .A2 (nx37296)) ;
    or03 ix24810 (.Y (nx24809), .A0 (nx37298), .A1 (nx37190), .A2 (nx37008)) ;
    or03 ix24817 (.Y (nx24816), .A0 (nx37002), .A1 (nx37190), .A2 (nx37298)) ;
    or03 ix24826 (.Y (nx24825), .A0 (nx36996), .A1 (nx37190), .A2 (nx37298)) ;
    or03 ix24831 (.Y (nx24830), .A0 (nx36990), .A1 (nx37190), .A2 (nx37298)) ;
    or03 ix24839 (.Y (nx24838), .A0 (nx36984), .A1 (nx37190), .A2 (nx37298)) ;
    or03 ix24846 (.Y (nx24845), .A0 (nx36978), .A1 (nx37190), .A2 (nx37300)) ;
    or03 ix24854 (.Y (nx24853), .A0 (nx36966), .A1 (nx37192), .A2 (nx37300)) ;
    or03 ix24860 (.Y (nx24859), .A0 (nx36972), .A1 (nx37192), .A2 (nx37300)) ;
    or03 ix24870 (.Y (nx24869), .A0 (nx36960), .A1 (nx37192), .A2 (nx37300)) ;
    or03 ix24875 (.Y (nx24874), .A0 (nx36954), .A1 (nx37192), .A2 (nx37300)) ;
    or03 ix24883 (.Y (nx24882), .A0 (nx36942), .A1 (nx37192), .A2 (nx37300)) ;
    or03 ix24888 (.Y (nx24887), .A0 (nx36948), .A1 (nx37192), .A2 (nx37300)) ;
    or03 ix24895 (.Y (nx24894), .A0 (nx36936), .A1 (nx37192), .A2 (nx37302)) ;
    or03 ix24901 (.Y (nx24900), .A0 (nx36930), .A1 (nx37194), .A2 (nx37302)) ;
    or03 ix24910 (.Y (nx24909), .A0 (nx36924), .A1 (nx37194), .A2 (nx37302)) ;
    or03 ix24915 (.Y (nx24914), .A0 (nx36916), .A1 (nx37194), .A2 (nx37302)) ;
    mux21 ix24922 (.Y (nx24921), .A0 (camera_module_algo_module_address_value_1)
          , .A1 (nx23005), .S0 (camera_module_algo_module_address_value_2)) ;
    ao32 ix753 (.Y (nx752), .A0 (nx22935), .A1 (nx22585), .A2 (nx22943), .B0 (
         camera_module_algo_module_address_value_0), .B1 (nx408)) ;
    mux21 ix17061 (.Y (nx17060), .A0 (nx35674), .A1 (nx24945), .S0 (nx37138)) ;
    mux21 ix24961 (.Y (nx24960), .A0 (nx14410), .A1 (nx14382), .S0 (nx37106)) ;
    mux21_ni ix14383 (.Y (nx14382), .A0 (nx14378), .A1 (nx14366), .S0 (nx37098)
             ) ;
    mux21_ni ix14367 (.Y (nx14366), .A0 (nvm_data_116), .A1 (nvm_data_124), .S0 (
             nx37160)) ;
    mux21_ni ix14379 (.Y (nx14378), .A0 (nvm_data_100), .A1 (nvm_data_108), .S0 (
             nx37160)) ;
    mux21_ni ix14411 (.Y (nx14410), .A0 (nx14406), .A1 (nx14394), .S0 (nx37098)
             ) ;
    mux21_ni ix14395 (.Y (nx14394), .A0 (nvm_data_84), .A1 (nvm_data_92), .S0 (
             nx37160)) ;
    mux21_ni ix14407 (.Y (nx14406), .A0 (nvm_data_68), .A1 (nvm_data_76), .S0 (
             nx37160)) ;
    mux21_ni ix14357 (.Y (nx14356), .A0 (nx14324), .A1 (nx14350), .S0 (nx37108)
             ) ;
    mux21_ni ix14351 (.Y (nx14350), .A0 (nx14346), .A1 (nx14334), .S0 (nx37100)
             ) ;
    mux21_ni ix14335 (.Y (nx14334), .A0 (nvm_data_52), .A1 (nvm_data_60), .S0 (
             nx37160)) ;
    mux21_ni ix14347 (.Y (nx14346), .A0 (nvm_data_36), .A1 (nvm_data_44), .S0 (
             nx37160)) ;
    mux21 ix24998 (.Y (nx24997), .A0 (nvm_data_20), .A1 (nvm_data_28), .S0 (
          nx37160)) ;
    mux21 ix11513 (.Y (nx11512), .A0 (nx35674), .A1 (nx26370), .S0 (nx37138)) ;
    mux21 ix26386 (.Y (nx26385), .A0 (nx8862), .A1 (nx8834), .S0 (nx37108)) ;
    mux21_ni ix8835 (.Y (nx8834), .A0 (nx8830), .A1 (nx8818), .S0 (nx37100)) ;
    mux21_ni ix8819 (.Y (nx8818), .A0 (nvm_data_114), .A1 (nvm_data_122), .S0 (
             nx37162)) ;
    mux21_ni ix8831 (.Y (nx8830), .A0 (nvm_data_98), .A1 (nvm_data_106), .S0 (
             nx37162)) ;
    mux21_ni ix8863 (.Y (nx8862), .A0 (nx8858), .A1 (nx8846), .S0 (nx37100)) ;
    mux21_ni ix8847 (.Y (nx8846), .A0 (nvm_data_82), .A1 (nvm_data_90), .S0 (
             nx37162)) ;
    mux21_ni ix8859 (.Y (nx8858), .A0 (nvm_data_66), .A1 (nvm_data_74), .S0 (
             nx37162)) ;
    mux21_ni ix8809 (.Y (nx8808), .A0 (nx8776), .A1 (nx8802), .S0 (nx37108)) ;
    mux21_ni ix8803 (.Y (nx8802), .A0 (nx8798), .A1 (nx8786), .S0 (nx37100)) ;
    mux21_ni ix8787 (.Y (nx8786), .A0 (nvm_data_50), .A1 (nvm_data_58), .S0 (
             nx37162)) ;
    mux21_ni ix8799 (.Y (nx8798), .A0 (nvm_data_34), .A1 (nvm_data_42), .S0 (
             nx37162)) ;
    mux21 ix26430 (.Y (nx26429), .A0 (nvm_data_18), .A1 (nvm_data_26), .S0 (
          nx37162)) ;
    mux21 ix5965 (.Y (nx5964), .A0 (nx35676), .A1 (nx27681), .S0 (nx37138)) ;
    mux21 ix27695 (.Y (nx27694), .A0 (nx1174), .A1 (nx1146), .S0 (nx37108)) ;
    mux21_ni ix1147 (.Y (nx1146), .A0 (nx1142), .A1 (nx1130), .S0 (nx37100)) ;
    mux21_ni ix1131 (.Y (nx1130), .A0 (nvm_data_112), .A1 (nvm_data_120), .S0 (
             nx37420)) ;
    mux21_ni ix1143 (.Y (nx1142), .A0 (nvm_data_96), .A1 (nvm_data_104), .S0 (
             nx37420)) ;
    mux21_ni ix1175 (.Y (nx1174), .A0 (nx1170), .A1 (nx1158), .S0 (nx37100)) ;
    mux21_ni ix1159 (.Y (nx1158), .A0 (nvm_data_80), .A1 (nvm_data_88), .S0 (
             nx37420)) ;
    mux21_ni ix1171 (.Y (nx1170), .A0 (nvm_data_64), .A1 (nvm_data_72), .S0 (
             nx37420)) ;
    mux21_ni ix1121 (.Y (nx1120), .A0 (nx1088), .A1 (nx1114), .S0 (nx37108)) ;
    mux21_ni ix1115 (.Y (nx1114), .A0 (nx1110), .A1 (nx1098), .S0 (nx37100)) ;
    mux21_ni ix1099 (.Y (nx1098), .A0 (nvm_data_48), .A1 (nvm_data_56), .S0 (
             nx37420)) ;
    mux21_ni ix1111 (.Y (nx1110), .A0 (nvm_data_32), .A1 (nvm_data_40), .S0 (
             nx37420)) ;
    mux21 ix27725 (.Y (nx27724), .A0 (nvm_data_16), .A1 (nvm_data_24), .S0 (
          nx37420)) ;
    xor2 ix28818 (.Y (nx28817), .A0 (nx29956), .A1 (nx28822)) ;
    mux21 ix8739 (.Y (nx8738), .A0 (nx35676), .A1 (nx28822), .S0 (nx37138)) ;
    mux21 ix28836 (.Y (nx28835), .A0 (nx6088), .A1 (nx6060), .S0 (nx37108)) ;
    mux21_ni ix6061 (.Y (nx6060), .A0 (nx6056), .A1 (nx6044), .S0 (nx37102)) ;
    mux21_ni ix6045 (.Y (nx6044), .A0 (nvm_data_113), .A1 (nvm_data_121), .S0 (
             nx37164)) ;
    mux21_ni ix6057 (.Y (nx6056), .A0 (nvm_data_97), .A1 (nvm_data_105), .S0 (
             nx37164)) ;
    mux21_ni ix6089 (.Y (nx6088), .A0 (nx6084), .A1 (nx6072), .S0 (nx37102)) ;
    mux21_ni ix6073 (.Y (nx6072), .A0 (nvm_data_81), .A1 (nvm_data_89), .S0 (
             nx37164)) ;
    mux21_ni ix6085 (.Y (nx6084), .A0 (nvm_data_65), .A1 (nvm_data_73), .S0 (
             nx37166)) ;
    mux21_ni ix6035 (.Y (nx6034), .A0 (nx6002), .A1 (nx6028), .S0 (nx37108)) ;
    mux21_ni ix6029 (.Y (nx6028), .A0 (nx6024), .A1 (nx6012), .S0 (nx37102)) ;
    mux21_ni ix6013 (.Y (nx6012), .A0 (nvm_data_49), .A1 (nvm_data_57), .S0 (
             nx37166)) ;
    mux21_ni ix6025 (.Y (nx6024), .A0 (nvm_data_33), .A1 (nvm_data_41), .S0 (
             nx37166)) ;
    mux21 ix28866 (.Y (nx28865), .A0 (nvm_data_17), .A1 (nvm_data_25), .S0 (
          nx37166)) ;
    xor2 ix29960 (.Y (nx29959), .A0 (nx31098), .A1 (nx29964)) ;
    mux21 ix14287 (.Y (nx14286), .A0 (nx35676), .A1 (nx29964), .S0 (nx37138)) ;
    mux21 ix29978 (.Y (nx29977), .A0 (nx11636), .A1 (nx11608), .S0 (nx37110)) ;
    mux21_ni ix11609 (.Y (nx11608), .A0 (nx11604), .A1 (nx11592), .S0 (nx37102)
             ) ;
    mux21_ni ix11593 (.Y (nx11592), .A0 (nvm_data_115), .A1 (nvm_data_123), .S0 (
             nx37166)) ;
    mux21_ni ix11605 (.Y (nx11604), .A0 (nvm_data_99), .A1 (nvm_data_107), .S0 (
             nx37166)) ;
    mux21_ni ix11637 (.Y (nx11636), .A0 (nx11632), .A1 (nx11620), .S0 (nx37102)
             ) ;
    mux21_ni ix11621 (.Y (nx11620), .A0 (nvm_data_83), .A1 (nvm_data_91), .S0 (
             nx37166)) ;
    mux21_ni ix11633 (.Y (nx11632), .A0 (nvm_data_67), .A1 (nvm_data_75), .S0 (
             nx37168)) ;
    mux21_ni ix11583 (.Y (nx11582), .A0 (nx11550), .A1 (nx11576), .S0 (nx37110)
             ) ;
    mux21_ni ix11577 (.Y (nx11576), .A0 (nx11572), .A1 (nx11560), .S0 (nx37102)
             ) ;
    mux21_ni ix11561 (.Y (nx11560), .A0 (nvm_data_51), .A1 (nvm_data_59), .S0 (
             nx37168)) ;
    mux21_ni ix11573 (.Y (nx11572), .A0 (nvm_data_35), .A1 (nvm_data_43), .S0 (
             nx37168)) ;
    mux21 ix30008 (.Y (nx30007), .A0 (nvm_data_19), .A1 (nvm_data_27), .S0 (
          nx37168)) ;
    xor2 ix31102 (.Y (nx31101), .A0 (nx32240), .A1 (nx31106)) ;
    mux21 ix19835 (.Y (nx19834), .A0 (nx35676), .A1 (nx31106), .S0 (nx37140)) ;
    mux21 ix31120 (.Y (nx31119), .A0 (nx17184), .A1 (nx17156), .S0 (nx37110)) ;
    mux21_ni ix17157 (.Y (nx17156), .A0 (nx17152), .A1 (nx17140), .S0 (nx37102)
             ) ;
    mux21_ni ix17141 (.Y (nx17140), .A0 (nvm_data_117), .A1 (nvm_data_125), .S0 (
             nx37168)) ;
    mux21_ni ix17153 (.Y (nx17152), .A0 (nvm_data_101), .A1 (nvm_data_109), .S0 (
             nx37168)) ;
    mux21_ni ix17185 (.Y (nx17184), .A0 (nx17180), .A1 (nx17168), .S0 (nx37104)
             ) ;
    mux21_ni ix17169 (.Y (nx17168), .A0 (nvm_data_85), .A1 (nvm_data_93), .S0 (
             nx37168)) ;
    mux21_ni ix17181 (.Y (nx17180), .A0 (nvm_data_69), .A1 (nvm_data_77), .S0 (
             nx37170)) ;
    mux21_ni ix17131 (.Y (nx17130), .A0 (nx17098), .A1 (nx17124), .S0 (nx37110)
             ) ;
    mux21_ni ix17125 (.Y (nx17124), .A0 (nx17120), .A1 (nx17108), .S0 (nx37104)
             ) ;
    mux21_ni ix17109 (.Y (nx17108), .A0 (nvm_data_53), .A1 (nvm_data_61), .S0 (
             nx37170)) ;
    mux21_ni ix17121 (.Y (nx17120), .A0 (nvm_data_37), .A1 (nvm_data_45), .S0 (
             nx37170)) ;
    mux21 ix31150 (.Y (nx31149), .A0 (nvm_data_21), .A1 (nvm_data_29), .S0 (
          nx37170)) ;
    xor2 ix32244 (.Y (nx32243), .A0 (nx33382), .A1 (nx32248)) ;
    mux21 ix25383 (.Y (nx25382), .A0 (nx35678), .A1 (nx32248), .S0 (nx37140)) ;
    mux21 ix32262 (.Y (nx32261), .A0 (nx22732), .A1 (nx22704), .S0 (nx37110)) ;
    mux21_ni ix22705 (.Y (nx22704), .A0 (nx22700), .A1 (nx22688), .S0 (nx37104)
             ) ;
    mux21_ni ix22689 (.Y (nx22688), .A0 (nvm_data_119), .A1 (nvm_data_127), .S0 (
             nx37170)) ;
    mux21_ni ix22701 (.Y (nx22700), .A0 (nvm_data_103), .A1 (nvm_data_111), .S0 (
             nx37170)) ;
    mux21_ni ix22733 (.Y (nx22732), .A0 (nx22728), .A1 (nx22716), .S0 (nx37104)
             ) ;
    mux21_ni ix22717 (.Y (nx22716), .A0 (nvm_data_87), .A1 (nvm_data_95), .S0 (
             nx37170)) ;
    mux21_ni ix22729 (.Y (nx22728), .A0 (nvm_data_71), .A1 (nvm_data_79), .S0 (
             nx35720)) ;
    mux21_ni ix22679 (.Y (nx22678), .A0 (nx22646), .A1 (nx22672), .S0 (nx37110)
             ) ;
    mux21_ni ix22673 (.Y (nx22672), .A0 (nx22668), .A1 (nx22656), .S0 (nx37104)
             ) ;
    mux21_ni ix22657 (.Y (nx22656), .A0 (nvm_data_55), .A1 (nvm_data_63), .S0 (
             nx35720)) ;
    mux21_ni ix22669 (.Y (nx22668), .A0 (nvm_data_39), .A1 (nvm_data_47), .S0 (
             nx35720)) ;
    mux21 ix32292 (.Y (nx32291), .A0 (nvm_data_23), .A1 (nvm_data_31), .S0 (
          nx35720)) ;
    xor2 ix26027 (.Y (nx26026), .A0 (nx25398), .A1 (nx37086)) ;
    xor2 ix33461 (.Y (nx33460), .A0 (nx22689), .A1 (nx37086)) ;
    xor2 ix26175 (.Y (nx26174), .A0 (nx25406), .A1 (nx37088)) ;
    xor2 ix33468 (.Y (nx33467), .A0 (nx22685), .A1 (nx37088)) ;
    xor2 ix26323 (.Y (nx26322), .A0 (nx25414), .A1 (nx37088)) ;
    xor2 ix33475 (.Y (nx33474), .A0 (nx22681), .A1 (nx37088)) ;
    nor03_2x ix693 (.Y (nx34150), .A0 (nx37084), .A1 (nx37416), .A2 (nx686)) ;
    mux21_ni ix22204 (.Y (nx22203), .A0 (
             camera_module_algo_module_current_cont_value_13), .A1 (nx26380), .S0 (
             nx37306)) ;
    mux21_ni ix26381 (.Y (nx26380), .A0 (
             camera_module_algo_module_Addout_value_13), .A1 (zero), .S0 (
             nx37074)) ;
    mux21_ni ix22194 (.Y (nx22193), .A0 (nx26366), .A1 (
             camera_module_algo_module_Addout_value_13), .S0 (nx37118)) ;
    mux21_ni ix26367 (.Y (nx26366), .A0 (zero), .A1 (nx26358), .S0 (nx37140)) ;
    mux21 ix22154 (.Y (nx22153), .A0 (nx33491), .A1 (nx33489), .S0 (nx37130)) ;
    mux21_ni ix22144 (.Y (nx22143), .A0 (
             camera_module_algo_module_current_cont_value_11), .A1 (nx26232), .S0 (
             nx37306)) ;
    mux21_ni ix26233 (.Y (nx26232), .A0 (
             camera_module_algo_module_Addout_value_11), .A1 (zero), .S0 (
             nx37074)) ;
    mux21_ni ix22134 (.Y (nx22133), .A0 (nx26218), .A1 (
             camera_module_algo_module_Addout_value_11), .S0 (nx37118)) ;
    mux21_ni ix26219 (.Y (nx26218), .A0 (zero), .A1 (nx26210), .S0 (nx37140)) ;
    mux21 ix22094 (.Y (nx22093), .A0 (nx33510), .A1 (nx33508), .S0 (nx37130)) ;
    mux21_ni ix22084 (.Y (nx22083), .A0 (
             camera_module_algo_module_current_cont_value_9), .A1 (nx26084), .S0 (
             nx37306)) ;
    mux21_ni ix26085 (.Y (nx26084), .A0 (
             camera_module_algo_module_Addout_value_9), .A1 (zero), .S0 (nx37074
             )) ;
    mux21_ni ix22074 (.Y (nx22073), .A0 (nx26070), .A1 (
             camera_module_algo_module_Addout_value_9), .S0 (nx37118)) ;
    mux21_ni ix26071 (.Y (nx26070), .A0 (zero), .A1 (nx26062), .S0 (nx37140)) ;
    mux21_ni ix22034 (.Y (nx22033), .A0 (nx25972), .A1 (
             camera_module_algo_module_diff_value_7), .S0 (nx37130)) ;
    mux21_ni ix25973 (.Y (nx25972), .A0 (zero), .A1 (nx25964), .S0 (nx37140)) ;
    mux21 ix25965 (.Y (nx25964), .A0 (nx33453), .A1 (nx33529), .S0 (nx37090)) ;
    mux21_ni ix22024 (.Y (nx22023), .A0 (
             camera_module_algo_module_current_cont_value_7), .A1 (nx25936), .S0 (
             nx37306)) ;
    mux21_ni ix25937 (.Y (nx25936), .A0 (
             camera_module_algo_module_Addout_value_7), .A1 (zero), .S0 (nx37074
             )) ;
    mux21_ni ix22014 (.Y (nx22013), .A0 (nx25922), .A1 (
             camera_module_algo_module_Addout_value_7), .S0 (nx37118)) ;
    mux21_ni ix25923 (.Y (nx25922), .A0 (zero), .A1 (nx25914), .S0 (nx37140)) ;
    mux21_ni ix21974 (.Y (nx21973), .A0 (nx25824), .A1 (
             camera_module_algo_module_diff_value_5), .S0 (nx37130)) ;
    mux21_ni ix25825 (.Y (nx25824), .A0 (zero), .A1 (nx25816), .S0 (nx37142)) ;
    mux21 ix25817 (.Y (nx25816), .A0 (nx33446), .A1 (nx33546), .S0 (nx37090)) ;
    mux21_ni ix21964 (.Y (nx21963), .A0 (
             camera_module_algo_module_current_cont_value_5), .A1 (nx25788), .S0 (
             nx37306)) ;
    mux21_ni ix25789 (.Y (nx25788), .A0 (
             camera_module_algo_module_Addout_value_5), .A1 (zero), .S0 (nx37370
             )) ;
    mux21_ni ix21954 (.Y (nx21953), .A0 (nx25774), .A1 (
             camera_module_algo_module_Addout_value_5), .S0 (nx37118)) ;
    mux21_ni ix25775 (.Y (nx25774), .A0 (zero), .A1 (nx25766), .S0 (nx37142)) ;
    mux21_ni ix21914 (.Y (nx21913), .A0 (nx25676), .A1 (
             camera_module_algo_module_diff_value_3), .S0 (nx37130)) ;
    mux21_ni ix25677 (.Y (nx25676), .A0 (zero), .A1 (nx25668), .S0 (nx37142)) ;
    mux21 ix25669 (.Y (nx25668), .A0 (nx33439), .A1 (nx33563), .S0 (nx37090)) ;
    mux21_ni ix21904 (.Y (nx21903), .A0 (
             camera_module_algo_module_current_cont_value_3), .A1 (nx25640), .S0 (
             nx37306)) ;
    mux21_ni ix25641 (.Y (nx25640), .A0 (
             camera_module_algo_module_Addout_value_3), .A1 (zero), .S0 (nx37370
             )) ;
    mux21_ni ix21894 (.Y (nx21893), .A0 (nx25626), .A1 (
             camera_module_algo_module_Addout_value_3), .S0 (nx37120)) ;
    mux21_ni ix25627 (.Y (nx25626), .A0 (zero), .A1 (nx25618), .S0 (nx37142)) ;
    mux21_ni ix21854 (.Y (nx21853), .A0 (nx25528), .A1 (
             camera_module_algo_module_diff_value_1), .S0 (nx37130)) ;
    mux21_ni ix25529 (.Y (nx25528), .A0 (zero), .A1 (nx25520), .S0 (nx37142)) ;
    mux21 ix25521 (.Y (nx25520), .A0 (nx33429), .A1 (nx33580), .S0 (nx37090)) ;
    mux21_ni ix21844 (.Y (nx21843), .A0 (
             camera_module_algo_module_current_cont_value_1), .A1 (nx25492), .S0 (
             nx37308)) ;
    mux21_ni ix25493 (.Y (nx25492), .A0 (
             camera_module_algo_module_Addout_value_1), .A1 (zero), .S0 (nx37370
             )) ;
    mux21_ni ix21834 (.Y (nx21833), .A0 (nx25478), .A1 (
             camera_module_algo_module_Addout_value_1), .S0 (nx37120)) ;
    mux21_ni ix25479 (.Y (nx25478), .A0 (zero), .A1 (nx25470), .S0 (nx37142)) ;
    xnor2 ix33592 (.Y (nx33591), .A0 (nx33609), .A1 (nx33615)) ;
    mux21_ni ix1244 (.Y (nx1243), .A0 (
             camera_module_algo_module_current_cont_value_0), .A1 (nx678), .S0 (
             nx37308)) ;
    mux21_ni ix679 (.Y (nx678), .A0 (camera_module_algo_module_Addout_value_0), 
             .A1 (zero), .S0 (nx37372)) ;
    mux21_ni ix1234 (.Y (nx1233), .A0 (nx664), .A1 (
             camera_module_algo_module_Addout_value_0), .S0 (nx37120)) ;
    mux21_ni ix665 (.Y (nx664), .A0 (zero), .A1 (nx656), .S0 (nx37142)) ;
    nor03_2x ix655 (.Y (nx34007), .A0 (nx37416), .A1 (
             camera_module_algo_module_modCU_current_state_5), .A2 (nx37070)) ;
    nand03 ix33602 (.Y (nx37070), .A0 (nx22993), .A1 (nx22979), .A2 (nx37072)) ;
    inv01 ix37071 (.Y (nx37072), .A (
          camera_module_algo_module_modCU_current_state_7)) ;
    nand04 ix33605 (.Y (nx36796), .A0 (nx37406), .A1 (nx37094), .A2 (nx22987), .A3 (
           nx33608)) ;
    mux21_ni ix21824 (.Y (nx21823), .A0 (nx25454), .A1 (
             camera_module_algo_module_diff_value_0), .S0 (nx37132)) ;
    mux21_ni ix25455 (.Y (nx25454), .A0 (zero), .A1 (nx25446), .S0 (nx37144)) ;
    mux21_ni ix25447 (.Y (nx25446), .A0 (nx25434), .A1 (nx25438), .S0 (nx37092)
             ) ;
    xor2 ix33617 (.Y (nx33616), .A0 (nx33619), .A1 (
         camera_module_algo_module_diff_value_1)) ;
    xnor2 ix33622 (.Y (nx33621), .A0 (nx33632), .A1 (nx33638)) ;
    mux21_ni ix21874 (.Y (nx21873), .A0 (
             camera_module_algo_module_current_cont_value_2), .A1 (nx25566), .S0 (
             nx37308)) ;
    mux21_ni ix25567 (.Y (nx25566), .A0 (
             camera_module_algo_module_Addout_value_2), .A1 (zero), .S0 (nx37372
             )) ;
    mux21_ni ix21864 (.Y (nx21863), .A0 (nx25552), .A1 (
             camera_module_algo_module_Addout_value_2), .S0 (nx37120)) ;
    mux21 ix25553 (.Y (nx25552), .A0 (nx35680), .A1 (nx33629), .S0 (nx37144)) ;
    mux21_ni ix21884 (.Y (nx21883), .A0 (nx25602), .A1 (
             camera_module_algo_module_diff_value_2), .S0 (nx37132)) ;
    mux21_ni ix25603 (.Y (nx25602), .A0 (zero), .A1 (nx25594), .S0 (nx37144)) ;
    mux21_ni ix25595 (.Y (nx25594), .A0 (nx25582), .A1 (nx25586), .S0 (nx37092)
             ) ;
    xor2 ix33640 (.Y (nx33639), .A0 (nx33642), .A1 (
         camera_module_algo_module_diff_value_3)) ;
    xnor2 ix33645 (.Y (nx33644), .A0 (nx33655), .A1 (nx33661)) ;
    mux21_ni ix21934 (.Y (nx21933), .A0 (
             camera_module_algo_module_current_cont_value_4), .A1 (nx25714), .S0 (
             nx37308)) ;
    mux21_ni ix25715 (.Y (nx25714), .A0 (
             camera_module_algo_module_Addout_value_4), .A1 (zero), .S0 (nx37372
             )) ;
    mux21_ni ix21924 (.Y (nx21923), .A0 (nx25700), .A1 (
             camera_module_algo_module_Addout_value_4), .S0 (nx37120)) ;
    mux21 ix25701 (.Y (nx25700), .A0 (nx35680), .A1 (nx33652), .S0 (nx37144)) ;
    mux21_ni ix21944 (.Y (nx21943), .A0 (nx25750), .A1 (
             camera_module_algo_module_diff_value_4), .S0 (nx37132)) ;
    mux21_ni ix25751 (.Y (nx25750), .A0 (zero), .A1 (nx25742), .S0 (nx37144)) ;
    mux21_ni ix25743 (.Y (nx25742), .A0 (nx25730), .A1 (nx25734), .S0 (nx37092)
             ) ;
    xor2 ix33663 (.Y (nx33662), .A0 (nx33665), .A1 (
         camera_module_algo_module_diff_value_5)) ;
    xnor2 ix33668 (.Y (nx33667), .A0 (nx33678), .A1 (nx33684)) ;
    mux21_ni ix21994 (.Y (nx21993), .A0 (
             camera_module_algo_module_current_cont_value_6), .A1 (nx25862), .S0 (
             nx37308)) ;
    mux21_ni ix25863 (.Y (nx25862), .A0 (
             camera_module_algo_module_Addout_value_6), .A1 (zero), .S0 (nx37372
             )) ;
    mux21_ni ix21984 (.Y (nx21983), .A0 (nx25848), .A1 (
             camera_module_algo_module_Addout_value_6), .S0 (nx37120)) ;
    mux21 ix25849 (.Y (nx25848), .A0 (nx35680), .A1 (nx33675), .S0 (nx37144)) ;
    mux21_ni ix22004 (.Y (nx22003), .A0 (nx25898), .A1 (
             camera_module_algo_module_diff_value_6), .S0 (nx37132)) ;
    mux21_ni ix25899 (.Y (nx25898), .A0 (zero), .A1 (nx25890), .S0 (nx37144)) ;
    mux21_ni ix25891 (.Y (nx25890), .A0 (nx25878), .A1 (nx25882), .S0 (nx37092)
             ) ;
    xor2 ix33686 (.Y (nx33685), .A0 (nx33688), .A1 (
         camera_module_algo_module_diff_value_7)) ;
    xnor2 ix33691 (.Y (nx33690), .A0 (nx33701), .A1 (nx33707)) ;
    mux21_ni ix22054 (.Y (nx22053), .A0 (
             camera_module_algo_module_current_cont_value_8), .A1 (nx26010), .S0 (
             nx37308)) ;
    mux21_ni ix26011 (.Y (nx26010), .A0 (
             camera_module_algo_module_Addout_value_8), .A1 (zero), .S0 (nx37074
             )) ;
    mux21_ni ix22044 (.Y (nx22043), .A0 (nx25996), .A1 (
             camera_module_algo_module_Addout_value_8), .S0 (nx37120)) ;
    mux21 ix25997 (.Y (nx25996), .A0 (nx35680), .A1 (nx33698), .S0 (nx35688)) ;
    mux21_ni ix22064 (.Y (nx22063), .A0 (nx26046), .A1 (
             camera_module_algo_module_diff_value_8), .S0 (nx37132)) ;
    mux21_ni ix26047 (.Y (nx26046), .A0 (zero), .A1 (nx26038), .S0 (nx35688)) ;
    mux21_ni ix26039 (.Y (nx26038), .A0 (nx26026), .A1 (nx26030), .S0 (nx37092)
             ) ;
    xnor2 ix33709 (.Y (nx33708), .A0 (nx33711), .A1 (nx33508)) ;
    xnor2 ix33714 (.Y (nx33713), .A0 (nx33724), .A1 (nx33727)) ;
    mux21_ni ix22114 (.Y (nx22113), .A0 (
             camera_module_algo_module_current_cont_value_10), .A1 (nx26158), .S0 (
             nx37308)) ;
    mux21_ni ix26159 (.Y (nx26158), .A0 (
             camera_module_algo_module_Addout_value_10), .A1 (zero), .S0 (
             nx37076)) ;
    mux21_ni ix22104 (.Y (nx22103), .A0 (nx26144), .A1 (
             camera_module_algo_module_Addout_value_10), .S0 (nx37122)) ;
    mux21 ix26145 (.Y (nx26144), .A0 (nx35680), .A1 (nx33721), .S0 (nx35688)) ;
    mux21 ix22124 (.Y (nx22123), .A0 (nx33729), .A1 (nx33727), .S0 (nx37132)) ;
    xnor2 ix33735 (.Y (nx33734), .A0 (nx33737), .A1 (nx33489)) ;
    xnor2 ix33740 (.Y (nx33739), .A0 (nx33750), .A1 (nx33753)) ;
    mux21_ni ix22174 (.Y (nx22173), .A0 (
             camera_module_algo_module_current_cont_value_12), .A1 (nx26306), .S0 (
             nx37310)) ;
    mux21_ni ix26307 (.Y (nx26306), .A0 (
             camera_module_algo_module_Addout_value_12), .A1 (zero), .S0 (
             nx37076)) ;
    mux21_ni ix22164 (.Y (nx22163), .A0 (nx26292), .A1 (
             camera_module_algo_module_Addout_value_12), .S0 (nx37122)) ;
    mux21 ix26293 (.Y (nx26292), .A0 (nx35682), .A1 (nx33747), .S0 (nx35688)) ;
    mux21 ix22184 (.Y (nx22183), .A0 (nx33755), .A1 (nx33753), .S0 (nx37132)) ;
    xnor2 ix33761 (.Y (nx33760), .A0 (nx33763), .A1 (nx22651)) ;
    xnor2 ix33766 (.Y (nx33765), .A0 (nx33776), .A1 (nx33779)) ;
    mux21_ni ix22234 (.Y (nx22233), .A0 (
             camera_module_algo_module_current_cont_value_14), .A1 (nx26454), .S0 (
             nx37310)) ;
    mux21_ni ix26455 (.Y (nx26454), .A0 (
             camera_module_algo_module_Addout_value_14), .A1 (zero), .S0 (
             nx37076)) ;
    mux21_ni ix22224 (.Y (nx22223), .A0 (nx26440), .A1 (
             camera_module_algo_module_Addout_value_14), .S0 (nx37122)) ;
    mux21 ix26441 (.Y (nx26440), .A0 (nx35682), .A1 (nx33773), .S0 (nx37146)) ;
    mux21 ix22244 (.Y (nx22243), .A0 (nx33781), .A1 (nx33779), .S0 (nx37134)) ;
    xor2 ix26471 (.Y (nx26470), .A0 (nx25422), .A1 (nx37088)) ;
    xnor2 ix33791 (.Y (nx33790), .A0 (nx33810), .A1 (nx33794)) ;
    mux21 ix22254 (.Y (nx22253), .A0 (nx33796), .A1 (nx33794), .S0 (nx37134)) ;
    xor2 ix33808 (.Y (nx33807), .A0 (nx22669), .A1 (nx37088)) ;
    mux21_ni ix22284 (.Y (nx22283), .A0 (
             camera_module_algo_module_prev_cont_value_15), .A1 (nx26580), .S0 (
             nx37076)) ;
    mux21_ni ix26581 (.Y (nx26580), .A0 (zero), .A1 (
             camera_module_algo_module_current_cont_value_15), .S0 (nx37146)) ;
    mux21_ni ix22294 (.Y (nx22293), .A0 (
             camera_module_algo_module_prev_cont_value_14), .A1 (nx26596), .S0 (
             nx37076)) ;
    mux21_ni ix26597 (.Y (nx26596), .A0 (zero), .A1 (
             camera_module_algo_module_current_cont_value_14), .S0 (nx37146)) ;
    xnor2 ix26605 (.Y (nx26604), .A0 (nx33776), .A1 (nx33818)) ;
    xnor2 ix33826 (.Y (nx33825), .A0 (nx33763), .A1 (
          camera_module_algo_module_prev_cont_value_13)) ;
    mux21_ni ix22304 (.Y (nx22303), .A0 (
             camera_module_algo_module_prev_cont_value_13), .A1 (nx26612), .S0 (
             nx37076)) ;
    mux21_ni ix26613 (.Y (nx26612), .A0 (zero), .A1 (
             camera_module_algo_module_current_cont_value_13), .S0 (nx37148)) ;
    mux21_ni ix22314 (.Y (nx22313), .A0 (
             camera_module_algo_module_prev_cont_value_12), .A1 (nx26628), .S0 (
             nx37076)) ;
    mux21_ni ix26629 (.Y (nx26628), .A0 (zero), .A1 (
             camera_module_algo_module_current_cont_value_12), .S0 (nx37148)) ;
    xnor2 ix26637 (.Y (nx26636), .A0 (nx33750), .A1 (nx33834)) ;
    xnor2 ix33842 (.Y (nx33841), .A0 (nx33737), .A1 (
          camera_module_algo_module_prev_cont_value_11)) ;
    mux21_ni ix22324 (.Y (nx22323), .A0 (
             camera_module_algo_module_prev_cont_value_11), .A1 (nx26644), .S0 (
             nx37078)) ;
    mux21_ni ix26645 (.Y (nx26644), .A0 (zero), .A1 (
             camera_module_algo_module_current_cont_value_11), .S0 (nx37148)) ;
    mux21_ni ix22334 (.Y (nx22333), .A0 (
             camera_module_algo_module_prev_cont_value_10), .A1 (nx26660), .S0 (
             nx37078)) ;
    mux21_ni ix26661 (.Y (nx26660), .A0 (zero), .A1 (
             camera_module_algo_module_current_cont_value_10), .S0 (nx37148)) ;
    xnor2 ix26669 (.Y (nx26668), .A0 (nx33724), .A1 (nx33850)) ;
    xnor2 ix33858 (.Y (nx33857), .A0 (nx33711), .A1 (
          camera_module_algo_module_prev_cont_value_9)) ;
    mux21_ni ix22344 (.Y (nx22343), .A0 (
             camera_module_algo_module_prev_cont_value_9), .A1 (nx26676), .S0 (
             nx37078)) ;
    mux21_ni ix26677 (.Y (nx26676), .A0 (zero), .A1 (
             camera_module_algo_module_current_cont_value_9), .S0 (nx37148)) ;
    mux21_ni ix22354 (.Y (nx22353), .A0 (
             camera_module_algo_module_prev_cont_value_8), .A1 (nx26692), .S0 (
             nx37078)) ;
    mux21_ni ix26693 (.Y (nx26692), .A0 (zero), .A1 (
             camera_module_algo_module_current_cont_value_8), .S0 (nx37148)) ;
    xnor2 ix26701 (.Y (nx26700), .A0 (nx33701), .A1 (nx33866)) ;
    xnor2 ix33874 (.Y (nx33873), .A0 (nx33688), .A1 (
          camera_module_algo_module_prev_cont_value_7)) ;
    mux21_ni ix22364 (.Y (nx22363), .A0 (
             camera_module_algo_module_prev_cont_value_7), .A1 (nx26708), .S0 (
             nx37078)) ;
    mux21_ni ix26709 (.Y (nx26708), .A0 (zero), .A1 (
             camera_module_algo_module_current_cont_value_7), .S0 (nx37148)) ;
    mux21_ni ix22374 (.Y (nx22373), .A0 (
             camera_module_algo_module_prev_cont_value_6), .A1 (nx26724), .S0 (
             nx37078)) ;
    mux21_ni ix26725 (.Y (nx26724), .A0 (zero), .A1 (
             camera_module_algo_module_current_cont_value_6), .S0 (nx37150)) ;
    xnor2 ix26733 (.Y (nx26732), .A0 (nx33678), .A1 (nx33882)) ;
    xnor2 ix33890 (.Y (nx33889), .A0 (nx33665), .A1 (
          camera_module_algo_module_prev_cont_value_5)) ;
    mux21_ni ix22384 (.Y (nx22383), .A0 (
             camera_module_algo_module_prev_cont_value_5), .A1 (nx26740), .S0 (
             nx37078)) ;
    mux21_ni ix26741 (.Y (nx26740), .A0 (zero), .A1 (
             camera_module_algo_module_current_cont_value_5), .S0 (nx37150)) ;
    mux21_ni ix22394 (.Y (nx22393), .A0 (
             camera_module_algo_module_prev_cont_value_4), .A1 (nx26756), .S0 (
             nx37080)) ;
    mux21_ni ix26757 (.Y (nx26756), .A0 (zero), .A1 (
             camera_module_algo_module_current_cont_value_4), .S0 (nx37150)) ;
    xnor2 ix26765 (.Y (nx26764), .A0 (nx33655), .A1 (nx33898)) ;
    xnor2 ix33906 (.Y (nx33905), .A0 (nx33642), .A1 (
          camera_module_algo_module_prev_cont_value_3)) ;
    mux21_ni ix22404 (.Y (nx22403), .A0 (
             camera_module_algo_module_prev_cont_value_3), .A1 (nx26772), .S0 (
             nx37080)) ;
    mux21_ni ix26773 (.Y (nx26772), .A0 (zero), .A1 (
             camera_module_algo_module_current_cont_value_3), .S0 (nx37150)) ;
    mux21_ni ix22414 (.Y (nx22413), .A0 (
             camera_module_algo_module_prev_cont_value_2), .A1 (nx26788), .S0 (
             nx37080)) ;
    mux21_ni ix26789 (.Y (nx26788), .A0 (zero), .A1 (
             camera_module_algo_module_current_cont_value_2), .S0 (nx37150)) ;
    xnor2 ix26797 (.Y (nx26796), .A0 (nx33632), .A1 (nx33914)) ;
    xnor2 ix33922 (.Y (nx33921), .A0 (nx33619), .A1 (
          camera_module_algo_module_prev_cont_value_1)) ;
    mux21_ni ix22424 (.Y (nx22423), .A0 (
             camera_module_algo_module_prev_cont_value_1), .A1 (nx26804), .S0 (
             nx37080)) ;
    mux21_ni ix26805 (.Y (nx26804), .A0 (zero), .A1 (
             camera_module_algo_module_current_cont_value_1), .S0 (nx37150)) ;
    mux21_ni ix22434 (.Y (nx22433), .A0 (
             camera_module_algo_module_prev_cont_value_0), .A1 (nx26820), .S0 (
             nx37080)) ;
    mux21_ni ix26821 (.Y (nx26820), .A0 (zero), .A1 (
             camera_module_algo_module_current_cont_value_0), .S0 (nx37150)) ;
    xnor2 ix26829 (.Y (nx26828), .A0 (nx33609), .A1 (nx33930)) ;
    mux21_ni ix22464 (.Y (nx22463), .A0 (
             camera_module_algo_module_current_cont_value_16), .A1 (nx27016), .S0 (
             nx37310)) ;
    mux21_ni ix27017 (.Y (nx27016), .A0 (
             camera_module_algo_module_Addout_value_16), .A1 (zero), .S0 (
             nx37080)) ;
    mux21_ni ix22454 (.Y (nx22453), .A0 (nx27002), .A1 (
             camera_module_algo_module_Addout_value_16), .S0 (nx37122)) ;
    mux21 ix27003 (.Y (nx27002), .A0 (nx35682), .A1 (nx33943), .S0 (nx35690)) ;
    mux21_ni ix22444 (.Y (nx22443), .A0 (nx26984), .A1 (
             camera_module_algo_module_diff_value_16), .S0 (nx37134)) ;
    xor2 ix33959 (.Y (nx33958), .A0 (zero), .A1 (nx37092)) ;
    nor02ii ix33962 (.Y (nx33961), .A0 (camera_module_algo_module_pixel_value_8)
            , .A1 (zero)) ;
    mux21_ni ix22474 (.Y (nx22473), .A0 (
             camera_module_algo_module_prev_cont_value_16), .A1 (nx27030), .S0 (
             nx37080)) ;
    mux21_ni ix27031 (.Y (nx27030), .A0 (zero), .A1 (
             camera_module_algo_module_current_cont_value_16), .S0 (nx35690)) ;
    or02 ix34004 (.Y (nx34003), .A0 (rst), .A1 (nx22601)) ;
    or02 ix34026 (.Y (nx20), .A0 (camera_module_ack_from_DMA), .A1 (rst)) ;
    and02 ix35705 (.Y (nx35706), .A0 (nx35688), .A1 (nx22601)) ;
    and02 ix35715 (.Y (nx35716), .A0 (nx37126), .A1 (nx37176)) ;
    and02 ix35797 (.Y (nx35798), .A0 (nx37406), .A1 (nx22979)) ;
    inv02 ix37073 (.Y (nx37074), .A (nx37406)) ;
    inv02 ix37075 (.Y (nx37076), .A (nx37406)) ;
    inv02 ix37077 (.Y (nx37078), .A (nx37406)) ;
    inv02 ix37079 (.Y (nx37080), .A (nx37114)) ;
    buf02 ix37081 (.Y (nx37082), .A (nx688)) ;
    buf02 ix37083 (.Y (nx37084), .A (nx688)) ;
    inv02 ix37085 (.Y (nx37086), .A (nx22677)) ;
    inv02 ix37087 (.Y (nx37088), .A (nx22677)) ;
    inv02 ix37089 (.Y (nx37090), .A (nx35700)) ;
    inv02 ix37091 (.Y (nx37092), .A (nx35700)) ;
    inv02 ix37093 (.Y (nx37094), .A (nx408)) ;
    inv02 ix37095 (.Y (nx37096), .A (nx34098)) ;
    inv02 ix37097 (.Y (nx37098), .A (nx34098)) ;
    inv02 ix37099 (.Y (nx37100), .A (nx34098)) ;
    inv02 ix37101 (.Y (nx37102), .A (nx34098)) ;
    inv02 ix37103 (.Y (nx37104), .A (nx34098)) ;
    inv02 ix37105 (.Y (nx37106), .A (nx34112)) ;
    inv02 ix37107 (.Y (nx37108), .A (nx34112)) ;
    inv02 ix37109 (.Y (nx37110), .A (nx34112)) ;
    inv02 ix37111 (.Y (nx37112), .A (nx404)) ;
    inv02 ix37113 (.Y (nx37114), .A (nx404)) ;
    inv01 ix37115 (.Y (nx37116), .A (nx34007)) ;
    inv02 ix37117 (.Y (nx37118), .A (nx37116)) ;
    inv02 ix37119 (.Y (nx37120), .A (nx37116)) ;
    inv02 ix37121 (.Y (nx37122), .A (nx37116)) ;
    inv02 ix37123 (.Y (nx37124), .A (camera_module_DMA_module_signals_1)) ;
    inv02 ix37125 (.Y (nx37126), .A (camera_module_DMA_module_signals_1)) ;
    inv01 ix37127 (.Y (nx37128), .A (nx34150)) ;
    inv02 ix37129 (.Y (nx37130), .A (nx37128)) ;
    inv02 ix37131 (.Y (nx37132), .A (nx37128)) ;
    inv02 ix37133 (.Y (nx37134), .A (nx37128)) ;
    inv02 ix37135 (.Y (nx37136), .A (nx37416)) ;
    inv02 ix37137 (.Y (nx37138), .A (nx37416)) ;
    inv02 ix37139 (.Y (nx37140), .A (nx37418)) ;
    inv02 ix37141 (.Y (nx37142), .A (nx37418)) ;
    inv02 ix37143 (.Y (nx37144), .A (nx37418)) ;
    inv02 ix37145 (.Y (nx37146), .A (nx37418)) ;
    inv02 ix37147 (.Y (nx37148), .A (nx37418)) ;
    inv02 ix37149 (.Y (nx37150), .A (nx37418)) ;
    buf02 ix37151 (.Y (nx37152), .A (nx35706)) ;
    buf02 ix37153 (.Y (nx37154), .A (nx35716)) ;
    inv02 ix37155 (.Y (nx37156), .A (nx37412)) ;
    inv02 ix37157 (.Y (nx37158), .A (nx37412)) ;
    inv02 ix37159 (.Y (nx37160), .A (nx37412)) ;
    inv02 ix37161 (.Y (nx37162), .A (nx37412)) ;
    inv02 ix37163 (.Y (nx37164), .A (nx37412)) ;
    inv02 ix37165 (.Y (nx37166), .A (nx37414)) ;
    inv02 ix37167 (.Y (nx37168), .A (nx37414)) ;
    inv02 ix37169 (.Y (nx37170), .A (nx37414)) ;
    inv02 ix37171 (.Y (nx37172), .A (nx37364)) ;
    inv02 ix37173 (.Y (nx37174), .A (nx37366)) ;
    inv02 ix37175 (.Y (nx37176), .A (nx37366)) ;
    inv02 ix37177 (.Y (nx37178), .A (nx37366)) ;
    inv02 ix37179 (.Y (nx37180), .A (nx37366)) ;
    inv02 ix37181 (.Y (nx37182), .A (nx37366)) ;
    inv02 ix37183 (.Y (nx37184), .A (nx37366)) ;
    inv02 ix37185 (.Y (nx37186), .A (nx37366)) ;
    inv02 ix37187 (.Y (nx37188), .A (nx37368)) ;
    inv02 ix37189 (.Y (nx37190), .A (nx37368)) ;
    inv02 ix37191 (.Y (nx37192), .A (nx36912)) ;
    inv02 ix37193 (.Y (nx37194), .A (nx36912)) ;
    inv02 ix37195 (.Y (nx37196), .A (nx436)) ;
    buf02 ix37197 (.Y (nx37198), .A (nx35798)) ;
    inv02 ix37199 (.Y (nx37200), .A (nx37012)) ;
    inv02 ix37201 (.Y (nx37202), .A (nx37006)) ;
    inv02 ix37203 (.Y (nx37204), .A (nx37000)) ;
    inv02 ix37205 (.Y (nx37206), .A (nx36994)) ;
    inv02 ix37207 (.Y (nx37208), .A (nx36988)) ;
    inv02 ix37209 (.Y (nx37210), .A (nx36982)) ;
    inv02 ix37211 (.Y (nx37212), .A (nx36970)) ;
    inv02 ix37213 (.Y (nx37214), .A (nx36976)) ;
    inv02 ix37215 (.Y (nx37216), .A (nx36964)) ;
    inv02 ix37217 (.Y (nx37218), .A (nx36958)) ;
    inv02 ix37219 (.Y (nx37220), .A (nx36946)) ;
    inv02 ix37221 (.Y (nx37222), .A (nx36952)) ;
    inv02 ix37223 (.Y (nx37224), .A (nx36940)) ;
    inv02 ix37225 (.Y (nx37226), .A (nx36934)) ;
    inv02 ix37227 (.Y (nx37228), .A (nx36928)) ;
    inv02 ix37229 (.Y (nx37230), .A (nx36920)) ;
    inv02 ix37231 (.Y (nx37232), .A (nx5650)) ;
    inv02 ix37233 (.Y (nx37234), .A (nx5650)) ;
    inv02 ix37235 (.Y (nx37236), .A (nx5358)) ;
    inv02 ix37237 (.Y (nx37238), .A (nx5358)) ;
    inv02 ix37239 (.Y (nx37240), .A (nx5064)) ;
    inv02 ix37241 (.Y (nx37242), .A (nx5064)) ;
    inv02 ix37243 (.Y (nx37244), .A (nx4772)) ;
    inv02 ix37245 (.Y (nx37246), .A (nx4772)) ;
    inv02 ix37247 (.Y (nx37248), .A (nx4474)) ;
    inv02 ix37249 (.Y (nx37250), .A (nx4474)) ;
    inv02 ix37251 (.Y (nx37252), .A (nx4182)) ;
    inv02 ix37253 (.Y (nx37254), .A (nx4182)) ;
    inv02 ix37255 (.Y (nx37256), .A (nx3888)) ;
    inv02 ix37257 (.Y (nx37258), .A (nx3888)) ;
    inv02 ix37259 (.Y (nx37260), .A (nx3596)) ;
    inv02 ix37261 (.Y (nx37262), .A (nx3596)) ;
    inv02 ix37263 (.Y (nx37264), .A (nx3294)) ;
    inv02 ix37265 (.Y (nx37266), .A (nx3294)) ;
    inv02 ix37267 (.Y (nx37268), .A (nx3002)) ;
    inv02 ix37269 (.Y (nx37270), .A (nx3002)) ;
    inv02 ix37271 (.Y (nx37272), .A (nx2708)) ;
    inv02 ix37273 (.Y (nx37274), .A (nx2708)) ;
    inv02 ix37275 (.Y (nx37276), .A (nx2416)) ;
    inv02 ix37277 (.Y (nx37278), .A (nx2416)) ;
    inv02 ix37279 (.Y (nx37280), .A (nx36506)) ;
    inv02 ix37281 (.Y (nx37282), .A (nx36506)) ;
    inv02 ix37283 (.Y (nx37284), .A (nx36506)) ;
    inv02 ix37285 (.Y (nx37286), .A (nx36580)) ;
    inv02 ix37287 (.Y (nx37288), .A (nx36580)) ;
    inv02 ix37289 (.Y (nx37290), .A (nx36580)) ;
    inv02 ix37291 (.Y (nx37292), .A (nx36654)) ;
    inv02 ix37293 (.Y (nx37294), .A (nx36654)) ;
    inv02 ix37295 (.Y (nx37296), .A (nx36654)) ;
    inv02 ix37297 (.Y (nx37298), .A (nx24811)) ;
    inv02 ix37299 (.Y (nx37300), .A (nx24811)) ;
    inv02 ix37301 (.Y (nx37302), .A (nx24811)) ;
    inv01 ix37303 (.Y (nx37304), .A (nx36796)) ;
    inv02 ix37305 (.Y (nx37306), .A (nx37304)) ;
    inv02 ix37307 (.Y (nx37308), .A (nx37304)) ;
    inv02 ix37309 (.Y (nx37310), .A (nx37304)) ;
    inv02 ix37311 (.Y (nx37312), .A (nx37422)) ;
    inv02 ix37313 (.Y (nx37314), .A (nx37422)) ;
    inv02 ix37315 (.Y (nx37316), .A (nx37422)) ;
    inv02 ix37317 (.Y (nx37318), .A (nx37422)) ;
    inv02 ix37319 (.Y (nx37320), .A (nx37422)) ;
    inv02 ix37321 (.Y (nx37322), .A (nx37422)) ;
    inv02 ix37323 (.Y (nx37324), .A (nx37424)) ;
    inv02 ix37325 (.Y (nx37326), .A (nx37424)) ;
    inv02 ix37327 (.Y (nx37328), .A (nx37424)) ;
    inv02 ix37329 (.Y (nx37330), .A (nx37424)) ;
    inv02 ix37331 (.Y (nx37332), .A (nx37424)) ;
    inv02 ix37333 (.Y (nx37334), .A (nx37424)) ;
    inv02 ix37335 (.Y (nx37336), .A (nx37424)) ;
    inv02 ix37337 (.Y (nx37338), .A (nx37426)) ;
    inv02 ix37339 (.Y (nx37340), .A (nx37426)) ;
    inv02 ix37341 (.Y (nx37342), .A (nx37426)) ;
    inv02 ix37343 (.Y (nx37344), .A (nx37426)) ;
    inv02 ix37345 (.Y (nx37346), .A (nx37426)) ;
    inv02 ix37347 (.Y (nx37348), .A (nx37426)) ;
    inv02 ix37349 (.Y (nx37350), .A (nx37426)) ;
    inv02 ix37351 (.Y (nx37352), .A (nx37428)) ;
    inv02 ix37353 (.Y (nx37354), .A (nx37428)) ;
    inv02 ix37355 (.Y (nx37356), .A (nx37428)) ;
    inv02 ix37357 (.Y (nx37358), .A (nx37428)) ;
    inv02 ix37359 (.Y (nx37360), .A (nx37428)) ;
    inv02 ix37361 (.Y (nx37362), .A (nx37428)) ;
    inv02 ix37363 (.Y (nx37364), .A (nx37428)) ;
    inv02 ix37365 (.Y (nx37366), .A (nx37430)) ;
    inv02 ix37367 (.Y (nx37368), .A (nx37430)) ;
    inv02 ix37369 (.Y (nx37370), .A (nx37112)) ;
    inv02 ix37371 (.Y (nx37372), .A (nx37112)) ;
    inv02 ix37373 (.Y (nx37374), .A (nx23298)) ;
    inv02 ix37375 (.Y (nx37376), .A (nx23290)) ;
    inv02 ix37377 (.Y (nx37378), .A (nx23279)) ;
    inv02 ix37379 (.Y (nx37380), .A (nx23267)) ;
    inv02 ix37381 (.Y (nx37382), .A (nx36208)) ;
    inv02 ix37383 (.Y (nx37384), .A (nx36248)) ;
    inv02 ix37385 (.Y (nx37386), .A (nx36168)) ;
    inv02 ix37387 (.Y (nx37388), .A (nx36128)) ;
    inv02 ix37389 (.Y (nx37390), .A (nx36048)) ;
    inv02 ix37391 (.Y (nx37392), .A (nx36088)) ;
    inv02 ix37393 (.Y (nx37394), .A (nx36008)) ;
    inv02 ix37395 (.Y (nx37396), .A (nx35968)) ;
    inv02 ix37397 (.Y (nx37398), .A (nx35928)) ;
    inv02 ix37399 (.Y (nx37400), .A (nx35888)) ;
    inv02 ix37401 (.Y (nx37402), .A (nx35848)) ;
    inv02 ix37403 (.Y (nx37404), .A (nx35808)) ;
    inv02 ix37405 (.Y (nx37406), .A (nx404)) ;
    inv02 ix37411 (.Y (nx37412), .A (nx35718)) ;
    inv02 ix37413 (.Y (nx37414), .A (nx35718)) ;
    inv02 ix37415 (.Y (nx37416), .A (nx35686)) ;
    inv02 ix37417 (.Y (nx37418), .A (nx35686)) ;
    inv02 ix37419 (.Y (nx37420), .A (camera_module_cache_address_from_DMA_0)) ;
    inv02 ix37421 (.Y (nx37422), .A (nx37436)) ;
    inv02 ix37423 (.Y (nx37424), .A (nx37438)) ;
    inv02 ix37425 (.Y (nx37426), .A (nx37438)) ;
    inv02 ix37427 (.Y (nx37428), .A (nx37438)) ;
    inv02 ix37429 (.Y (nx37430), .A (nx37438)) ;
    inv02 ix37435 (.Y (nx37436), .A (nx37028)) ;
    inv02 ix37437 (.Y (nx37438), .A (nx37028)) ;
endmodule

